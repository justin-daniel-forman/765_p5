`timescale 1ns/100ps
// VERILOG TESTBENCH// TB_justin_s9234_scan.v
// Input file: justin_s9234_scan.vectors.stil
// Converted from stil to Verilog TestBench
//
// Module "modulename"
// 925 vectors in file
// 1 clock signals present
// 38 input signals present (not including clocks)
// 40 output signals preset
//
// CLOCKS: CK
// INPUTS: TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23
// OUTPUTS: SO_TDI, g2584, g3222, g3600, g4307, g4321, g4422, g4809, g5137, g5468, g5469, g5692, g6282, g6284, g6360, g6362, g6364, g6366, g6368, g6370, g6372, g6374, g6728, g1290, g4121, g4108, g4106, g4103, g1293, g4099, g4102, g4109, g4100, g4112, g4105, g4101, g4110, g4104, g4107, g4098


module TB_modulename();
	wire SO_TDI, g2584, g3222, g3600, g4307, g4321, g4422, g4809, g5137, g5468, g5469, g5692, g6282, g6284, g6360, g6362, g6364, g6366, g6368, g6370, g6372, g6374, g6728, g1290, g4121, g4108, g4106, g4103, g1293, g4099, g4102, g4109, g4100, g4112, g4105, g4101, g4110, g4104, g4107, g4098;	//output signals
	reg CK, TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23;	//input signals

	//Insert correct wiring below
	modulename TOP (CLOCKS, INPUTS, OUTPUTS);

	initial begin
		CK = 1'b0;
		//Test vector 1
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'bZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		#5;
		CK = 1'b0;
		//Test vector 2
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b00ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 3
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b110ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 4
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b110ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 5
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 6
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 7
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 8
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 9
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 10
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b110ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 11
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b110ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 12
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 13
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 14
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b110ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 15
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 16
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 17
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 18
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 19
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 20
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 21
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 22
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 23
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 24
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 25
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 26
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 27
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 28
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 29
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 30
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 31
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 32
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 33
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 34
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 35
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 36
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 37
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 38
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 39
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 40
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 41
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 42
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 43
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 44
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 45
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 46
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 47
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 48
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 49
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 50
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 51
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 52
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 53
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 54
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 55
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 56
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 57
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 58
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 59
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 60
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 61
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 62
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 63
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 64
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 65
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 66
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 67
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 68
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 69
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 70
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 71
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 72
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 73
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 74
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 75
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 76
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 77
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 78
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 79
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 80
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 81
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 82
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 83
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 84
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 85
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 86
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 87
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 88
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 89
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 90
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 91
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 92
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 93
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 94
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 95
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 96
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 97
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 98
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 99
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 100
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 101
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 102
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 103
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 104
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 105
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 106
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 107
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 108
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 109
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 110
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 111
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 112
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 113
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 114
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 115
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 116
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 117
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 118
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 119
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 120
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 121
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 122
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 123
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 124
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 125
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 126
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 127
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 128
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 129
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 130
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 131
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 132
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 133
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 134
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 135
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 136
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 137
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 138
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 139
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 140
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 141
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 142
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 143
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 144
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 145
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 146
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 147
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 148
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 149
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 150
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 151
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 152
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 153
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 154
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 155
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 156
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 157
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 158
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 159
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 160
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 161
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 162
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 163
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 164
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 165
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 166
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 167
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 168
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 169
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 170
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 171
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 172
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 173
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 174
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 175
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 176
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 177
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 178
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 179
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 180
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 181
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 182
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 183
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 184
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 185
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 186
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 187
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 188
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 189
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 190
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 191
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 192
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 193
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 194
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 195
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 196
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 197
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 198
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 199
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 200
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 201
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 202
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 203
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 204
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 205
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 206
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 207
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 208
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 209
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 210
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 211
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 212
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 213
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 214
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 215
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 216
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 217
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 218
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 219
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 220
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 221
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 222
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 223
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 224
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 225
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 226
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 227
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 228
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b01Z110110000001101011001000110101101010;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 229
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b110ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 230
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b110ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 231
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 232
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 233
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b00ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 234
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b110ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 235
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b110ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 236
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 237
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 238
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 239
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 240
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 241
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b110ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 242
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b110ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 243
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 244
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 245
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b110ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 246
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 247
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 248
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 249
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 250
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 251
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 252
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 253
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 254
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 255
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 256
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 257
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 258
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 259
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 260
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 261
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 262
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 263
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 264
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 265
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 266
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 267
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 268
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 269
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 270
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 271
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 272
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 273
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 274
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 275
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 276
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 277
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 278
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 279
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 280
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 281
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 282
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 283
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 284
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 285
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 286
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 287
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 288
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 289
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 290
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 291
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 292
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 293
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 294
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 295
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 296
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 297
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 298
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 299
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 300
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 301
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 302
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 303
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 304
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 305
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 306
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 307
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 308
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 309
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 310
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 311
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 312
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 313
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 314
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 315
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 316
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 317
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 318
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 319
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 320
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 321
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 322
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 323
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 324
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 325
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 326
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 327
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 328
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 329
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 330
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 331
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 332
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 333
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 334
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 335
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 336
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 337
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 338
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 339
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 340
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 341
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 342
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 343
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 344
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 345
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 346
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 347
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 348
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 349
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 350
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 351
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 352
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 353
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 354
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 355
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 356
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 357
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 358
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 359
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 360
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 361
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 362
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 363
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 364
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 365
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 366
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 367
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 368
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 369
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 370
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 371
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 372
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 373
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 374
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 375
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 376
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 377
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 378
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 379
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 380
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 381
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 382
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 383
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 384
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 385
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 386
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 387
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 388
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 389
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 390
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 391
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 392
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 393
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 394
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 395
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 396
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 397
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 398
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 399
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 400
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 401
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 402
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 403
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 404
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 405
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 406
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 407
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 408
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 409
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 410
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 411
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 412
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 413
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 414
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 415
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 416
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 417
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 418
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 419
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 420
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 421
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 422
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 423
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 424
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 425
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 426
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 427
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 428
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 429
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 430
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 431
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 432
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 433
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 434
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 435
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 436
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 437
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 438
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 439
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 440
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 441
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 442
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 443
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 444
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 445
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 446
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 447
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 448
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 449
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 450
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 451
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 452
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 453
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 454
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 455
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 456
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 457
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 458
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 459
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b01Z101000100111011110111110110000001110;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 460
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b110ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 461
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b110ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 462
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 463
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 464
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b00ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 465
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b110ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 466
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b110ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 467
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 468
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 469
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 470
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 471
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 472
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b110ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 473
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b110ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 474
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 475
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 476
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b110ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 477
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 478
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 479
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 480
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 481
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 482
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 483
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 484
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 485
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 486
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 487
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 488
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 489
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 490
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 491
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 492
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 493
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 494
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 495
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 496
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 497
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 498
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 499
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 500
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 501
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 502
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 503
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 504
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 505
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 506
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 507
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 508
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 509
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 510
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 511
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 512
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 513
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 514
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 515
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 516
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 517
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 518
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 519
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 520
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 521
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 522
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 523
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 524
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 525
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 526
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 527
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 528
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 529
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 530
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 531
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 532
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 533
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 534
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 535
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 536
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 537
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 538
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 539
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 540
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 541
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 542
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 543
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 544
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 545
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 546
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 547
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 548
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 549
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 550
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 551
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 552
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 553
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 554
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 555
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 556
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 557
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 558
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 559
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 560
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 561
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 562
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 563
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 564
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 565
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 566
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 567
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 568
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 569
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 570
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 571
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 572
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 573
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 574
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 575
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 576
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 577
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 578
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 579
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 580
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 581
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 582
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 583
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 584
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 585
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 586
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 587
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 588
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 589
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 590
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 591
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 592
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 593
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 594
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 595
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 596
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 597
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 598
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 599
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 600
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 601
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 602
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 603
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 604
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 605
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 606
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 607
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 608
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 609
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 610
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 611
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 612
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 613
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 614
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 615
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 616
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 617
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 618
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 619
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 620
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 621
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 622
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 623
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 624
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 625
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 626
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 627
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 628
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 629
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 630
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 631
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 632
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 633
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 634
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 635
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 636
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 637
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 638
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 639
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 640
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 641
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 642
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 643
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 644
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 645
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 646
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 647
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 648
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 649
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 650
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 651
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 652
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 653
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 654
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 655
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 656
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 657
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 658
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 659
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 660
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 661
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 662
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 663
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 664
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 665
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 666
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 667
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 668
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 669
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 670
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 671
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 672
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 673
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 674
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 675
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 676
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 677
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 678
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 679
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 680
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 681
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 682
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 683
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 684
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 685
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 686
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 687
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 688
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 689
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 690
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b01Z000001111000101000010010110111101000;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 691
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b110ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 692
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b110ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 693
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 694
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 695
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b00ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 696
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b110ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 697
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b110ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 698
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 699
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 700
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 701
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 702
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 703
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b110ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 704
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b110ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 705
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 706
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 707
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b110ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 708
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 709
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 710
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 711
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 712
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 713
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 714
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 715
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 716
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 717
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 718
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 719
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 720
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 721
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 722
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 723
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 724
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 725
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 726
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 727
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 728
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 729
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 730
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 731
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 732
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 733
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 734
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 735
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 736
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 737
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 738
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 739
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 740
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 741
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 742
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 743
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 744
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 745
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 746
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 747
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 748
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 749
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 750
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 751
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 752
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 753
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 754
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 755
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 756
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 757
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 758
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 759
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 760
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 761
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 762
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 763
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 764
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 765
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 766
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 767
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 768
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 769
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 770
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 771
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 772
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 773
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 774
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 775
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 776
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 777
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 778
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 779
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 780
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 781
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 782
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 783
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 784
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 785
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 786
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 787
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 788
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 789
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 790
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 791
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 792
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 793
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 794
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 795
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 796
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 797
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 798
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 799
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 800
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 801
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 802
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 803
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 804
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 805
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 806
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 807
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 808
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 809
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 810
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 811
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 812
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 813
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 814
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 815
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 816
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 817
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 818
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 819
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 820
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 821
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 822
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 823
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 824
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 825
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 826
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 827
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 828
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 829
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 830
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 831
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 832
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 833
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 834
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 835
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 836
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 837
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 838
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 839
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 840
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 841
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 842
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 843
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 844
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 845
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 846
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 847
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 848
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 849
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 850
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 851
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 852
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 853
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 854
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 855
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 856
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 857
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 858
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 859
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 860
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 861
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 862
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 863
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 864
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 865
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 866
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 867
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 868
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 869
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 870
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 871
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 872
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 873
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 874
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 875
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 876
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 877
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 878
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 879
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 880
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 881
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 882
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 883
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 884
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 885
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 886
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 887
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 888
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 889
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 890
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 891
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 892
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 893
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 894
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 895
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 896
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 897
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 898
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 899
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 900
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 901
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 902
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 903
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 904
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 905
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 906
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 907
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 908
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 909
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 910
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 911
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 912
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 913
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 914
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 915
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 916
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 917
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 918
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 919
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b011ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 920
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 921
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b01ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 922
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b110ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 923
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b110ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 924
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
		CK = 1'b0;
		//Test vector 925
		{TMS, TRST, SI_TDI, g89, g94, g98, g102, g107, g301, g306, g310, g314, g319, g557, g558, g559, g560, g561, g562, g563, g564, g705, g639, g567, g45, g42, g39, g702, g32, g38, g46, g36, g47, g40, g37, g41, g22, g44, g23} = 39'b010ZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZZ;
		#5;
		CK = 1'b1;
		#5;
	end
endmodule
