// s9234 with its DFFs replaced with scan flip flops

module s9234_inscan(CK,g102,g107,g1290,g1293,g22,g23,g2584,g301,g306,g310,g314,g319,g32,
  g3222,g36,g3600,g37,g38,g39,g40,g4098,g4099,g41,g4100,g4101,g4102,g4103,
  g4104,g4105,g4106,g4107,g4108,g4109,g4110,g4112,g4121,g42,g4307,g4321,g44,
  g4422,g45,g46,g47,g4809,g5137,g5468,g5469,g557,g558,g559,g560,g561,g562,g563,
  g564,g567,g5692,g6282,g6284,g6360,g6362,g6364,g6366,g6368,g6370,g6372,g6374,
  g639,g6728,g702,g705,g89,g94,g98,clockdr,updatedr,shiftdr,TDI_ISR,TDO_ISR,int_hold,bistsel);

input CK,g89,g94,g98,g102,g107,g301,g306,g310,g314,g319,g557,g558,g559,g560,g561,
  g562,g563,g564,g705,g639,g567,g45,g42,g39,g702,g32,g38,g46,g36,g47,g40,g37,
  g41,g22,g44,g23,clockdr,updatedr,shiftdr,TDI_ISR,int_hold,bistsel;

output g2584,g3222,g3600,g4307,g4321,g4422,g4809,g5137,g5468,g5469,g5692,g6282,
  g6284,g6360,g6362,g6364,g6366,g6368,g6370,g6372,g6374,g6728,g1290,g4121,
  g4108,g4106,g4103,g1293,g4099,g4102,g4109,g4100,g4112,g4105,g4101,g4110,
  g4104,g4107,g4098,TDO_ISR;

  wire g678,g4130,g332,g6823,g123,g6940,g207,g6102,g695,g4147,g461,g4841,g18,
    g6725,g292,g3232,g331,g4119,g689,g4141,g24,g6726,g465,g6507,g84,g6590,g291,
    g3231,g676,g5330,g622,g5147,g117,g4839,g278,g6105,g128,g5138,g598,g4122,
    g554,g6827,g496,g6745,g179,g6405,g48,g6729,g590,g6595,g551,g6826,g682,
    g4134,g11,g6599,g606,g4857,g188,g6406,g646,g5148,g327,g4117,g361,g6582,
    g289,g3229,g398,g5700,g684,g4136,g619,g4858,g208,g5876,g248,g3239,g390,
    g5698,g625,g5328,g681,g4133,g437,g4847,g276,g5877,g3,g6597,g323,g4120,g224,
    g3235,g685,g4137,g43,g6407,g157,g5470,g282,g6841,g697,g4149,g206,g6101,
    g449,g4844,g118,g4113,g528,g6504,g284,g3224,g426,g4855,g634,g4424,g669,
    g5582,g520,g6502,g281,g6107,g175,g5472,g15,g6602,g631,g5581,g69,g6587,g693,
    g4145,g337,g2585,g457,g4842,g486,g2586,g471,g1291,g328,g4118,g285,g3225,
    g418,g4853,g402,g4849,g297,g6512,g212,g3233,g410,g4851,g430,g4856,g33,
    g6854,g662,g1831,g453,g4843,g269,g6510,g574,g6591,g441,g4846,g664,g1288,
    g349,g5478,g211,g6840,g586,g6594,g571,g5580,g29,g6853,g326,g4840,g698,
    g4150,g654,g5490,g293,g6511,g690,g4142,g445,g4845,g374,g5694,g6,g6722,g687,
    g4139,g357,g5480,g386,g5697,g504,g6498,g665,g4126,g166,g5471,g541,g6505,
    g74,g6588,g338,g5475,g696,g4148,g516,g6501,g536,g6506,g683,g4135,g353,
    g5479,g545,g6824,g254,g3240,g341,g5476,g290,g3230,g2,g6721,g287,g3227,g336,
    g6925,g345,g5477,g628,g5489,g679,g4131,g28,g6727,g688,g4140,g283,g6842,
    g613,g4423,g10,g6723,g14,g6724,g680,g4132,g143,g6401,g672,g5491,g667,g4127,
    g366,g6278,g279,g6106,g492,g6744,g170,g6404,g686,g4138,g288,g3228,g638,
    g1289,g602,g4123,g642,g4658,g280,g5878,g663,g4125,g610,g4124,g148,g5874,
    g209,g6103,g675,g1294,g478,g1292,g122,g4115,g54,g6584,g594,g6596,g286,
    g3226,g489,g2587,g616,g4657,g79,g6589,g218,g3234,g242,g3238,g578,g6592,
    g184,g5473,g119,g4114,g668,g6800,g139,g5141,g422,g4854,g210,g6839,g394,
    g5699,g230,g3236,g25,g6601,g204,g5875,g658,g4425,g650,g5329,g378,g5695,
    g508,g6499,g548,g6825,g370,g5693,g406,g4850,g236,g3237,g500,g6497,g205,
    g6100,g197,g6509,g666,g4128,g114,g4116,g524,g6503,g260,g3241,g111,g6277,
    g131,g5139,g7,g6598,g19,g6600,g677,g4129,g582,g6593,g485,g6801,g699,g4426,
    g193,g5474,g135,g5140,g382,g5696,g414,g4852,g434,g4848,g266,g4659,g49,
    g6583,g152,g6402,g692,g4144,g277,g6104,g127,g6941,g161,g6403,g512,g6500,
    g532,g6508,g64,g6586,g694,g4146,g691,g4143,g1,g6720,g59,g6585,I8854,g6696,
    I2272,I9125,g6855,I6783,g4822,I4424,g2097,g6895,I9152,g1835,I2919,I3040,
    g1770,g6837,g6822,I7466,g5624,I4809,g2974,g3537,I4757,g5457,g5304,g6062,
    g5824,g4040,I5343,I6001,g4162,g5549,g5331,I4477,g3063,g3612,I7055,g5318,
    g2892,g1982,I5264,g3638,I2225,I5451,g4323,g4086,g908,I1932,I5933,g4346,
    I8252,g6294,I2473,g971,I7333,g5386,I8812,g6688,g1674,g985,I3528,g1422,
    I8958,g6774,I5050,g3246,I4501,I2324,g1209,g2945,I4133,g5121,I6775,g1997,
    g1398,g3128,I4375,I8005,g6110,g1541,g1094,g5670,g5527,g2738,g2327,I9047,
    g4528,I6096,g2244,I3379,g6192,g5946,g2709,I3864,g1332,I2349,g4530,I6102,
    g1680,g1011,g2078,g1345,I2215,I3010,g1504,g5813,I7612,I7509,g5587,I5379,
    g3940,g3800,g3388,g2907,g1914,I9085,g2035,I3144,g2959,g1861,I9236,g4010,
    g3601,I2287,g927,I4273,g2197,I8270,g6300,g5740,I7501,I5777,g3807,g2876,
    g1943,g873,I6525,I5882,g3871,g2656,I3800,I8473,g6485,I2199,g900,I1927,
    g6708,I8834,I2399,g729,I3278,g1695,g6520,I8476,g940,I6677,g4757,g3902,
    g3575,g5687,g5567,g2915,g1931,g847,I3235,g1807,I3343,g1623,g6431,I8295,
    g709,g6812,I8984,I6576,g4700,g749,I1847,g3090,I4331,I9107,g2214,I3349,
    g4618,g4246,g6376,g6267,I5511,I6349,g4569,g4343,g4011,I5674,g4003,I8177,
    g6173,g2110,g1381,I3134,g1336,I8229,I3334,g1330,I7197,g5431,g4566,g4198,
    I7397,g5561,I4534,g2858,g1714,g1110,I4961,g3597,g2663,g2308,g3456,g2640,
    I6801,g922,I1947,g4693,I6283,I5484,g5570,g5392,g5860,g5634,g4334,g3733,
    I3804,g2575,I2207,I5153,g3330,g3355,g3100,g5645,g5537,g6733,I8891,g5691,
    g5568,g4804,g4473,g6838,I4414,g2090,g6610,I8696,g2877,g2434,I4903,g3223,
    g6796,I4288,I3313,g1337,g5879,g5770,g3463,g2682,I4513,g2765,I2578,g5358,
    I7012,I3202,g1812,I5421,g1076,I2115,g6069,g5791,I7817,g5924,g6540,g6474,
    I6352,g4564,I1865,g4202,I5622,I6867,g5082,g3876,I7349,I8144,g6182,g1175,
    g1375,I2411,g3118,I4366,g3318,I4593,g2464,I3596,g3872,g3312,g4494,I6004,
    I2870,g1161,g4518,I6066,g2215,g5615,I7372,g4567,I6139,I4382,g2265,I3776,
    g2044,g3057,I4282,I5600,g3821,I3593,g1295,I2825,g1143,g1285,g852,g3457,
    g2653,g5174,g5099,I6386,g4462,I3965,g2268,I8488,g6426,g6849,I9074,I6599,
    g4823,I2408,g719,g3834,I5027,g2295,g1578,g1384,I2420,g1339,I2370,g5545,
    I6170,I9128,g6864,g6898,I9161,g1838,g1595,g6900,I9167,g2194,I3331,g6797,
    I8961,g2394,I3537,I3050,g1439,I3641,g1491,I2943,g1715,I5736,g4022,I8450,
    I6280,g4430,g4933,I6625,g5420,I7086,g4521,I6075,g1672,I7058,g5281,I2887,
    g1123,I2122,g1477,g952,I4495,I2228,g5794,I7593,g1643,I2608,g3022,I4437,
    g2108,g2705,I3858,g3813,g3258,I8650,g6529,g1647,g2242,I3373,g1205,I2033,
    I5871,g3744,g774,I1859,g6819,I8994,g6694,I8800,g4379,I5848,g5905,g5852,
    g3519,g2740,I7856,g5994,g921,g1551,g1742,I2756,I4752,g2859,g6488,g6367,
    g2254,I3391,I8594,g6446,g2814,I4023,g4289,I5746,I6247,I6756,g4775,g6701,
    I8821,I8972,g6795,I3271,g1748,I2845,g1193,g5300,I6952,g2350,I3502,I8806,
    g6686,I3611,g1771,I2137,I8943,I2337,I2913,g1792,g1754,I2773,g6886,g2409,
    g1815,g894,I1917,g1273,g839,I5424,g3725,I6403,g4492,g6314,I8044,g4799,
    g4485,I9155,g6882,g2836,g2509,g2212,I6763,g4780,g3860,I5081,g2967,I4166,
    I9008,g5440,g5266,g3710,g3029,I5523,g3840,g843,g1543,g1006,I5478,g6408,
    g6283,g4153,I5545,I6359,g6136,g2822,I4031,g6706,I8913,g6743,I2692,g1037,
    g946,g1729,I2731,I5551,g4059,g4802,I6470,g3962,I5214,I2154,I4189,g2159,
    I5499,g3847,g5151,I6819,g3158,I4398,g6806,I8978,I4706,I7637,g5530,I7270,
    g6878,I5926,g2921,g1950,g6065,g5784,I6315,g4446,I4371,g2555,g6887,I4429,
    g2102,g6122,I7838,g6465,I8329,g6322,I8056,g1660,g1946,I3053,g6230,g6040,
    g5010,I6646,g4511,I6045,I6874,g4861,g2895,g1894,g6033,g2837,g2512,I2979,
    g1263,g5884,g5864,I8342,I2218,g1513,g878,I2312,g897,I3714,g1852,I4297,
    I8255,g6292,I8815,g6689,I5998,I1868,I7608,g5605,I5862,g3863,g1679,g1378,
    I2414,g4714,I6324,I2293,g5278,I6937,g3284,g3019,I4684,g2687,I8497,g6481,
    I4516,I6537,g4711,g3545,g3085,g2788,I3983,g6137,I7859,g5667,g5524,g6891,
    I9140,I2907,g1335,I2358,g3380,g2831,I4791,g6337,I8089,I4309,g2525,I2828,
    g3832,I5023,I2269,g5566,I7318,g3853,I5068,I3736,g2460,I6612,g4660,I7161,
    g5465,I7361,g2842,I4050,g1805,I2854,I6417,g4617,I3623,g4262,I5713,I7051,
    g5219,I2221,g3559,g2603,g4736,I6366,g2485,I3614,I7451,g5597,I2703,g1189,
    I8267,g6297,g4623,g1947,I3056,I5885,g3746,I7999,I7146,g5231,I6330,g4560,
    I7346,g5531,I3871,g2145,g6305,g4375,I5840,g4871,I8761,g6563,g3204,I4441,
    g4722,I6346,g710,I4498,g2686,g829,g5113,I6753,g1632,g760,I2067,I4347,I8828,
    g6661,I8872,I8411,g1653,I2630,I3782,I8727,g6536,g2031,I3140,I5436,g3729,
    g2252,I3385,g5908,g5753,g2958,I7472,g5626,g2176,I3319,I2716,g1115,I5831,
    g3842,g1160,I5182,g3271,g5518,I7258,g5418,I5382,g3952,g2405,I3543,I2848,
    g1917,I3016,g2829,g2491,I3946,I7116,g5299,I4019,g1841,I5923,I6090,g4393,
    I4362,I3672,g1656,g3040,I4255,I3077,I6485,g5593,I7355,g3440,I4678,g3969,
    I5233,g6312,I8040,I4452,g2117,I4173,I8217,g895,I6456,g4633,g4523,I6081,
    g1233,I2231,I6649,g4643,g4293,g5264,g4943,I9158,g1054,g5160,g2796,I3999,
    I6355,g2473,I3605,I3099,g1519,I8576,g6436,I2805,I8866,I3304,g1740,I4486,
    g3093,g5521,I7261,I3499,g1450,I8716,g6518,g1725,g1113,I7596,I8875,g3875,
    I5106,g2324,I3478,I4504,g2726,I2119,g5450,g5292,I5037,g3705,g5996,I5394,
    I8644,g4499,I6015,I2352,I6063,g4381,g6746,I8916,I2867,I8699,g6573,g2177,
    I3322,g5179,g5379,I7035,I2893,g1236,I7646,I3044,g1257,I2196,g3839,I5040,
    g6932,I9217,g4273,I5728,g5658,g5512,g6624,I8730,I6118,g4406,I6318,g4447,
    g2276,g2849,g2577,I3572,g1787,I2835,I5442,g3731,g2670,I6057,I8524,g6496,
    g6526,g1461,I6989,g5307,I2614,g1675,g1101,I2125,g3343,g3571,I2821,g1221,
    g4712,g6576,g6487,I6549,g4699,I8258,g6293,I8818,g6690,I3534,g2245,I3382,
    I3729,g2436,I3961,I5454,g3874,g2291,I3434,g5997,g5854,g4534,I6114,I3927,
    I5532,g3861,g1684,I2668,g6699,g1639,g815,g1338,I2367,g1963,I3074,I8186,
    g6179,I6321,g4559,I4226,g1109,g1791,I8975,g6791,g2256,g889,I2306,g896,
    g3792,g4745,g2819,g2467,g4014,I5316,I8426,g6424,I5412,g4034,I6253,g4608,
    g2088,g2923,g1969,g2408,I8614,g6537,I3513,g2488,I3617,g1759,I2782,g2701,
    I3855,I7190,g5432,g6691,g6524,I6740,g4781,g4513,I6051,g6794,g5596,g1957,
    I3068,I3352,g6119,I7829,I2904,g1256,g6319,I8051,g1049,g5901,g2886,g1966,
    I6552,g4702,I4059,g1878,g4036,I5337,g3094,I4337,I4459,g2134,I8544,g6453,
    g4679,I6269,g6352,I8110,g6818,I8991,g6577,I3288,g1710,g3567,g3074,g1284,
    I5487,I7704,g5723,g848,g5092,g4753,g1498,I2479,I2763,g2870,g2296,I3022,
    g1426,I4261,g1857,I2391,g4382,I5857,g3776,g3466,g6893,I9146,g1833,I3422,
    g1641,g5574,g5407,I3749,g2484,g3593,g2997,g6211,g5992,g2650,I3794,g5714,
    I7475,g932,I8061,g6113,g4805,I5328,g1584,g743,g4111,I8665,g1539,I5109,
    I3546,I2159,I6570,g4719,g2136,g1395,I4664,g2924,I8027,g6237,I4246,g2336,
    I3488,I7336,g716,I1832,I3560,g1673,g736,I1841,g4770,g2768,g2367,I8174,
    g2594,I3723,g4798,I6464,g6325,g6821,g6785,g4188,g2806,g2446,I3632,g3450,
    I4688,I3037,g1769,g6939,I9230,g1052,I3653,g1305,I3102,I2315,g1222,I2811,
    g6083,g5809,g2887,g1858,I2047,g6544,I6607,g4632,g4281,g5889,g5742,I7164,
    g2934,g2004,g2230,I3355,g4437,I5948,I5388,g4302,g4068,I5865,g3743,I7814,
    g4579,g4206,g4869,g4662,g6306,I8030,I3752,g5375,I7029,I8107,I6337,g1730,
    g1114,g3289,g3034,I2485,g3777,I6587,g4803,I8159,g6167,I6111,g4404,g3835,
    I5030,I6311,g4444,I8223,g2096,I3212,I9143,g3882,I5119,g1070,g2550,I3665,
    I6615,g3042,I4671,g2928,I2880,g2845,g2565,g1897,I2992,g6622,I8724,I2537,
    I5896,g3879,g2195,g4265,I5716,g2891,g1884,g2913,g1925,I6795,I3364,g1648,
    g5384,g5220,I9134,g6904,I9179,g4786,I6448,g3799,g6514,I8462,g4364,I5825,
    I8447,g6410,I3770,I5019,I2417,I7683,g5702,I9044,g3541,g2643,I2982,g1678,
    I2658,I6414,I2234,g1331,I2346,g4296,I5753,I2128,I3553,I6020,g4176,g3332,
    g3079,I7167,I6420,g6695,I8803,I2330,g1122,g3209,I6507,g4644,g4532,I6108,
    g1682,I9113,I1856,g3802,g2481,I3608,g5627,g931,g2692,I3840,I4217,g2163,
    I3215,I4066,g2582,g5551,I7295,g5686,I3886,I6737,g2497,I3626,I5385,I6956,
    g2154,g1755,I2776,g4189,I5597,g6792,g4706,I6308,g6416,I8243,g6286,I8417,
    g6420,g3901,I6630,g5774,I3675,g6522,I8482,g6115,g1045,I3281,g1761,I7039,
    g5309,I7484,g5630,g1173,I2185,I4455,g2118,I8629,g5273,I6930,g2040,I2476,
    I1853,g2783,I3979,g2112,I3240,g1283,g853,g2312,I3462,g1369,I2405,I6750,
    g4771,g6654,I8758,g3714,g3041,I7583,I3684,g1733,I5006,g3604,g6684,g1059,
    I2552,g2001,I3112,I5406,g3976,g5572,g5399,I3109,I3791,g2293,g1567,g6880,
    I8653,I5496,g1535,g1088,g4639,I8527,g5543,I3808,g2125,I7276,g3881,I2355,
    g1177,I5409,g4309,g4074,g2828,g2830,g2494,g2727,g4808,I2964,g821,I1880,
    g6612,I8702,g5534,g5729,I7494,I6666,g4740,g6875,g1415,g1246,g4707,g6417,
    I8261,I7404,g5541,g3076,I8512,g6441,g3889,I6528,g4815,g1664,I2643,I2237,
    g6234,g6057,I3575,g5885,g5865,g6328,I8066,g1203,I5445,g6542,I8538,g6330,
    I8070,g1721,I2721,I5091,g3242,g6109,g2932,g1998,I8456,g5903,I3833,g2266,
    I2318,g4715,I6327,I1924,I8966,I5169,I6410,I5376,g3500,g2647,g4498,I6012,
    I2057,g1502,I5059,g3259,I5920,g4228,I2457,g1253,I3584,I5868,g3864,I2989,
    I2193,g5436,g3384,g2834,g1940,I3047,g2576,I3687,g2866,g1905,g5135,g2716,
    g3838,I7906,g5912,I3268,I3019,g3424,g5382,I7042,I5793,g3803,I3419,g1287,
    g6902,I9173,I6143,g4237,I6343,g4458,g846,g1671,g5805,I7604,I5415,g3723,
    I3452,I5562,g5022,g1030,I8279,g6307,I4492,g6490,g6371,I2321,g898,I9002,
    g3477,g6166,I7892,I8162,I6334,g4454,g2241,I3370,g1564,g5916,I3086,I8503,
    I8843,g6658,g6649,I8745,I6555,g4703,g1741,I2753,I6792,g5097,g3104,I4351,
    g1318,g2524,I3647,g2644,I3788,g6698,g1638,g754,I6621,g2119,g1391,I5502,
    g1108,I2134,I3025,g5437,I7119,g4385,I3425,g1274,I9092,g2109,g2818,g2867,
    g1908,g1883,g1797,g5579,I7478,g5628,g5150,I7517,g2893,g1985,g5752,I8232,
    g6332,g5917,I6567,I3678,g1690,g2975,I4176,g1631,I2967,I8165,g1048,I5430,
    g3727,g2599,g5042,I6672,g1711,I2712,I3635,g6652,I8752,g5442,g5270,g1055,
    I2570,I2860,I5475,I4743,I3105,g2170,I3301,g2370,I3522,I5913,g6193,g5957,
    g1333,I3255,I8552,g6455,g1774,I2817,g4766,I6406,I5397,g1846,I2940,g5054,
    g4816,g4801,g4487,g6834,I5991,I7110,g5291,g3534,I5910,g3750,I3755,g5296,
    I6946,I8687,g6568,I6933,g5124,g2544,I3662,I8662,I5609,g3893,I4474,g3052,
    g1176,g3014,g6121,I7835,I7002,g5308,g766,g3885,I5124,g4226,g4050,g2106,
    g2306,g1743,g1320,g2790,g2413,g6232,g6048,I5217,g3673,I8570,g6433,I8860,
    I4480,g3073,g1994,I2275,g909,g6938,I9227,I5466,g3787,g4173,I5577,I8710,
    g6517,g2461,I7590,I3602,I3007,g2756,g2353,g2622,I3764,I3059,I3578,g1484,
    I3868,g5888,g5731,g838,g6519,I6289,g4433,I9024,g6803,I5448,g3960,I3767,
    g5787,g5685,g2904,g1991,g6552,g6606,I8684,I3581,I5333,g3491,I2284,g4718,
    g4767,g4601,I3261,g1783,g1847,g3207,I5774,I9077,g6845,I8659,g6523,g4535,
    I4976,g1685,I2671,I8506,g6483,g2841,g2541,g4582,g4210,I4229,g2391,I8626,
    I2029,g964,g791,g2695,I3843,g2637,I3779,g4227,g5439,g3798,I9104,g5063,
    I3284,g6570,I5692,I6132,g4219,g6525,I8491,g6710,I8840,I5418,I6680,g4713,
    g4721,I2588,g2416,I3556,g3095,I4340,g3037,I4252,g845,I2204,I5493,I8180,
    g6176,I4220,g2164,I7966,I8591,g6448,g2315,I3465,g5866,g6879,g6607,I6558,
    g4705,g4502,g5049,I6685,g6836,I1958,I1942,g3719,g3053,I8438,g5575,g5411,
    I8420,g6422,I3388,g1324,g2874,g1849,g3752,I4935,g3932,I3028,I5594,g4388,
    g3724,I3428,g1825,I2973,g1687,I7254,g5458,g5922,I3247,g6615,I8707,I7150,
    g5355,I4327,g4428,g3786,g5584,g5539,g5896,I2653,I3826,g3364,g3114,I8515,
    g6492,g4192,g3054,I4279,g4002,I4303,g2612,I8300,g6299,I8002,g2243,I3376,
    g3770,I9014,g6820,I3638,g1772,I5723,g3942,g4741,I6371,I8641,g5052,I6692,
    g6832,I9021,g4910,I2648,g980,g2234,I3367,I9082,g1890,g1359,I3883,g2574,
    I4240,g2165,g2330,g1777,g4609,I6182,I8441,g4308,I2050,g1734,I3758,g2041,
    g5086,g4732,g6142,g951,I8969,g2800,g2430,g5730,I7497,g2554,I3669,g4758,
    I6382,I2839,I3861,g1834,g6905,I9182,I3711,g1848,I4986,g2213,I3346,g5897,
    g5025,g4814,g6515,g5425,I7091,I2172,I2278,g917,I7796,I4681,g2947,g1480,
    g2902,g1899,g6697,I2143,I2343,g4222,I5481,g3297,g3046,I3206,I6546,I2334,
    I6809,g5051,I5743,I6995,I5890,g3878,I3509,g3963,g3791,I8884,g6704,I5505,
    g1688,I2688,g4752,I6434,I2961,I6231,g4350,g4509,I6039,g5087,I9095,g5801,
    I7600,g2155,I3274,I9208,g6922,g4640,I3093,g965,I3493,I3816,g2580,g1326,
    I8235,I6099,g4398,I8282,g6309,g3049,I4270,g6528,I8500,g1760,I2785,g4493,
    g6351,I1850,g834,I8988,g6787,g6530,I4777,g5045,I8693,g6655,g5445,g5274,
    I4799,I8548,g6454,I7193,g3498,g2634,I5854,g2619,I3761,I8555,g6456,I3519,
    g2872,g1922,g1608,g1220,I6292,I8240,I9164,g6885,g4397,I9233,g1192,I7640,
    g5773,I7073,g6884,I9119,I2593,g5059,I6697,g5920,I7692,I9038,g2457,I3587,
    g5578,I6444,g4503,g4655,g1423,I2442,g923,g3740,I7176,g1588,g798,I8113,
    g6147,I7342,I2182,I3830,g3162,I4402,g5261,I6918,I4294,I6543,g6618,g1665,
    g5926,g2158,g6143,I7865,g4562,g6235,g2598,I3726,g1327,I2521,g1063,g5415,
    I7081,g3452,g2625,I7996,I5400,g6566,I8582,I8494,g6428,I6534,I8518,g6494,
    g1681,g4723,I8567,g6432,g6134,I7852,g5664,g5352,g2232,I3361,g6548,I6927,
    g3086,I2724,g2253,I2179,g3486,g2869,g2813,I2379,g1696,I2700,I6885,g4872,
    g4497,g3504,g2675,g1732,I2738,I5116,I3909,g1001,I3441,I7069,g3070,I8264,
    g6296,g6621,I8721,I7469,g5625,g3897,g3251,g3263,g1472,g1043,I5977,g4319,
    I8521,g6495,I6036,g4370,I2611,g893,g6412,g1739,g1116,I3531,g1593,g3967,
    g4249,I8470,g6567,I8585,g6533,g4460,g996,I2041,g3331,I3890,g4772,g5247,
    g4900,g4531,I6105,I5633,g3768,I8878,I2663,I3505,I8647,g3766,I4955,g1533,
    g5564,I5103,I3650,g3801,g3487,I3013,I5696,g2691,g2317,I6798,g5741,g5602,
    I2802,g1204,I3474,g5638,g6160,I5508,g3867,g6933,I9220,I5944,g4356,g2962,
    g2008,g6521,I8479,I9098,I5472,g3846,I8981,g6793,g2506,I3080,I8674,g1820,
    I5043,g3247,I6495,g4607,g1936,g1756,I6437,g4501,g3173,I4410,g4399,I6302,
    g4440,I8997,g6790,g1117,I8541,g6452,g1317,g2608,I6579,g5993,g3557,I3569,
    g1789,g2111,g2275,g5466,I8332,I7701,g5720,g3369,I4646,I8153,g6185,g3007,
    g2615,I9101,I2864,g5571,g5395,g5861,g5636,g3868,g2174,g3459,g2664,I1877,
    g1775,g5448,g835,g5711,g6835,I9028,g1581,g910,I6042,g4374,g1060,g2284,
    I3431,I6786,g4824,g1460,g3793,g6611,g2591,I3720,g3015,I2749,I6054,g4194,
    g5538,I6296,g4436,g2602,I2623,I5460,g5509,I7251,g4400,I5899,g1937,g6541,
    I8535,I9185,g6877,I8600,g6451,g2931,g1988,g4760,I8074,g5067,g1190,I2175,
    g6353,g5873,g2905,g4167,I8910,g6802,g2628,g1156,g2515,g5493,I7065,g5256,
    g5077,I6706,g4731,g4220,I5644,I5177,I4276,I3161,g1270,g5381,I4667,I9131,
    g6901,I9170,g3771,I8623,g3216,g1824,g5552,I8453,g6457,I2424,I1844,g862,
    g2973,I4170,g1954,I3065,g3030,I4243,g1250,I5739,g1363,g1837,I5463,g5950,
    g1053,g1738,I8668,g6574,g6484,g2440,g3564,g2618,g6714,g6670,I5520,I5668,
    g3828,g4284,I8285,g6310,g3732,I5391,g6580,g6491,g6032,g5631,g5536,g3108,
    g6876,I6362,I4354,g3308,g3060,I6759,g4778,g2875,I6377,g4508,I8809,g6687,
    g6623,g6076,g5797,g6889,g5751,I7506,I3316,g1344,g3589,I7481,g5629,I3034,
    g2410,I3550,g1627,g2777,g6375,I8189,g2884,I2044,g3084,g2839,g2535,I5084,
    I7960,g5925,g899,g6651,I8749,g3448,g4565,g4195,I3681,g1821,I5053,g3455,
    g6285,g2172,I3307,g6937,I5568,g4533,g2667,I3811,g1683,g1017,g2343,g5168,
    g6339,I8093,g3196,I4433,g4914,I5002,I5630,I7267,I5157,g3454,I9035,I9203,
    g6921,g1731,I3258,g1735,I2745,I8273,g6301,g6809,g5890,g1782,g1935,I6452,
    g4629,I5929,g4152,g1661,g6252,g6231,g6044,g5011,I8444,g6421,g3067,g784,
    I1838,I7077,I8485,g861,I2946,g1587,g2792,I2584,I5433,I2281,I5626,g3914,
    I4334,g1646,I2617,g5869,g4191,g1084,I7808,g854,g1039,I2449,g6778,I6425,
    g5573,g5403,I5056,g4619,I2831,g2518,I3644,g1583,g1702,g1107,I2382,I8414,
    g6418,I8946,g1919,I2916,g2776,g2378,g4784,g1276,g2283,I3294,g1720,g3852,
    g6572,I4762,g2862,g5532,I6635,g2264,I3405,g6712,g6676,g851,I6766,g4783,
    I6087,g4392,g6543,I6305,g4441,g2360,g1793,g2933,I4123,I2620,g4190,I5526,
    g3848,g4157,I8335,g6308,I8831,g6665,g6931,g1546,I2873,I2037,g6534,I8881,
    g3605,I4802,I5603,g2996,I3942,g1503,I5439,g3730,g6742,g6560,g2179,I3328,
    g6014,I9122,g4704,g6414,I5702,g3845,I4258,g5383,I7045,g4903,g5303,g6903,
    I9176,g3441,g2835,g1407,g4250,g6513,I8459,g913,g4613,I5952,g4367,g4810,
    I6488,g2882,g1854,I7352,g5533,g3075,g872,g6036,I8632,I2364,g6531,I2808,
    g3772,I6582,g4765,I6689,g2981,I8579,g6438,I8869,I4489,g3458,g865,I2296,
    g3890,I4192,g4170,I3659,I4471,I7170,g5435,I8276,g4929,g2744,I1935,g2802,
    g2437,g949,I8564,I5320,g4626,g4270,g1340,I2373,g3480,g2986,g6653,I8755,
    I7802,I7061,I7187,g5387,g6579,g5116,I5987,g4224,g5316,I6976,I2635,g5434,
    g2864,g1887,I6430,g855,g4894,g4813,g1249,g4620,I5252,I2791,I7514,g5590,
    I2309,I2140,I8888,I3691,g5210,g6786,I6564,I8171,g6170,I8429,g6425,I7358,
    g6164,I8156,g6233,g6052,I2707,g4292,I7695,g2968,I5078,I2890,g4526,g3859,
    I7107,g5277,I5907,g3883,g1762,g2889,g1975,g4403,g4603,g6532,g4443,I5517,
    I9041,g4439,g5117,g6553,I5876,g3870,g2175,g2871,I2604,g3183,I4420,g2722,
    I4462,g2135,I8309,g6304,g1556,g3779,I8246,g3023,g1928,I3031,I7811,g5921,
    I7698,g1064,g6888,I2998,I6048,g4376,I7339,g4276,I5731,I4249,I3004,I1825,
    g4561,g2838,g1747,g3451,I2162,g1563,I9011,g2809,g1586,g4527,I6093,I2290,
    g4647,g3346,I4623,I5236,g2672,g2231,I3358,g4764,I6400,g5995,g6844,I7173,
    I3785,I6780,g4825,g1394,g1206,I6023,I2735,I2728,g1232,g1557,g4046,I5556,
    g2104,g1372,g2099,g1366,I4519,I2385,g6707,g1471,I2464,g4320,I3906,g4394,
    g6189,g3043,I4264,g3748,I6816,g5111,I3516,g2754,g2347,g4242,g1254,g1814,
    g6575,g6486,g4516,I6060,g6715,g6673,g4716,g5250,g6604,I8678,g1038,I6397,
    g1773,I2814,I2131,I7104,g4299,I5756,g6833,g6535,g5453,g2712,g2320,g6711,
    g4016,I8620,g6539,I8531,g6896,g1836,I2922,g5423,g6116,g6461,I8897,g1918,
    I3244,I7490,g5583,I4980,g3546,g5853,I4324,g2961,I5071,I3340,g1282,I5705,
    g6162,I8150,g6419,I6723,g4761,g2927,g1979,g4360,g6930,g2885,g5535,g6565,
    I2445,g2660,g2946,g938,g4435,g4517,g5717,I3656,I4794,I2491,g2903,g1902,
    I8635,g6363,I2169,g942,g6730,g3775,I8432,g3922,I7463,g5622,g6385,g6271,
    g6881,I9110,g3980,g2036,g1764,g706,I6441,g4624,g4915,g4669,g2178,I3325,
    g2679,I3823,g6070,I3525,I4285,I3310,g1640,g6897,I2925,g6561,g3460,I8226,
    I4510,g2753,g6890,g5452,I4291,g5894,g2805,g2443,I1938,g1788,g2422,I6772,
    g4788,g6480,I4312,I6531,g4402,g4017,I1862,I2240,g4615,g837,g5661,I1835,
    I3590,g1781,I7686,g5705,g1842,g1612,g1219,g6427,g6087,I6942,I8767,g6619,
    g6365,g3501,I3222,g1790,g6447,I6244,g6439,I2958,I9116,g6298,g5084,g4727,
    I5654,I3797,I6992,g2346,I5837,g3850,g2433,I2388,I6573,I3563,g6290,I2601,
    g2752,g6373,I8183,g3363,g3110,g5919,I7689,I2428,g4563,I2190,I3408,g3453,
    g6369,g2042,I3155,I5249,g6578,g6489,I6540,I3291,g1286,g2364,g2233,I5612,
    g1911,g5136,g3912,g3505,I2741,I8940,g6783,I2910,g1645,I3071,g5647,I3705,
    g2316,I3471,I2638,g844,g5546,g5388,g3857,I4465,g6015,g5857,g6415,I6126,
    g4240,I5686,I2883,I8671,I7707,g6239,g2103,I2327,I5708,I8857,I5640,g5120,
    g6429,g2706,I3773,I2165,I2212,g2888,g1972,g5565,I4195,g2173,g2029,g2171,
    g1934,g2787,g2956,g4151,I8638,I3819,I3836,g1832,g1806,I7587,g4769,g4606,
    I2949,g3778,g6188,I6949,g4185,g1898,I2995,g3782,g6562,g6114,g5892,g4451,
    I8290,I4306,g4229,I7284,g4614,g6564,I5324,I7832,g5943,I5469,g1953,g3267,
    I4321,g1819,I2877,g2957,g6685,I2952,I6072,g6609,I7113,I8034,I3062,g1776,
    g2449,I3620,g6450,g2865,g6883,g4837,I8509,g6437,g2604,I4267,g2098,g4251,
    g945,g6466,g5915,I7679,g4622,I8467,g6789,g6291,I2150,g6165,g6571,I8597,
    g5110,I5699,g5310,I3298,g1650,I2627,I3485,g3527,g809,I1874,g849,I5606,
    I5879,I2361,g3970,g1594,g6538,g6469,I3083,I2857,I7643,I3708,g2086,I3198,
    g2728,I4468,g2583,g3320,g6067,g5788,g1275,g6467,g1322,g4520,g1328,g4431,
    I5938,g4252,g1321,g3906,g2470,g3789,g5064,g2025,g6493,g5899,g4790,I5843,
    g4405,I4964,g1550,g4380,g4286,I4198,g3299,g5563,g4911,I3733,g6700,g1891,
    I2986,g5237,g5083,g3892,g2678,I3225,g1813,g6442,g4225,g2766,g2361,g2087,
    g1352,g2105,I7143,g5323,g2801,I4003,g5089,I5065,g714,I3540,g1670,g4980,
    g4678,g2748,I3923,g1823,g3478,g1142,g2755,g2169,g5242,g5085,I8168,I8863,
    g1255,I5033,I7799,g6817,g3728,g3082,I4315,g3482,g2713,g6444,g1692,I2696,
    g6605,I8681,g1726,g2091,g1355,g1960,g5295,g3751,g2061,g2007,g1411,I6250,
    g4514,g2059,g1402,g2920,g2157,g6118,g2767,I4358,I4821,I3090,g1112,g1267,
    g4510,g1319,g5918,g3002,I8573,g6435,I4483,I5514,I8713,I4507,g1329,I2340,
    I3694,g1811,I2788,g857,g5872,g2581,I2760,g3866,I8907,I9137,g1830,I7264,
    I8435,g6411,g6734,I8894,g1703,g4215,I5637,I2779,g6074,g3064,g3785,g1624,
    I2581,g5895,g4314,g4080,g6080,g1075,I8603,I4391,g6713,g6679,g1644,g6569,
    g2030,I3137,I5490,I4223,I8220,g4768,g2826,g1699,g4386,g2861,g4806,I8423,
    g6423,g5050,g1724,I8588,g6443,I4522,g1174,g842,g4434,g3083,g4322,I3232,
    g2609,g4687,g6527,g6108,I7153,g2883,I6084,g4391,g4182,I3096,I3496,g715,
    g5708,g1119,g2066,g1341,g3150,g1315,I8103,I3395,I3337,g4496,I6008,g1577,
    g4550,g3773,I4537,g5958,g5818,I2147,g6608,I8690,I5615,g830,g3769,g3622,
    g2827,g3856,g3836,g3212,g1853,g2333,g6287,g3844,g4807,I5223,I6561,I2596,
    g6161,g856,g6361,I8147,g2196,g2803,g4159,I6986,g5230,g6051,g804,I1871,
    g2538,g1325,I3481,g6242,g4248,g4692,I7805,I3599,g4726,g4154,I5548,g1636,
    g3921,g3512,g5540,g1106,g6732,I2842,I5893,g3747,I2460,g3462,g2381,I6789,
    g6043,I7871,g6097,I3001,g4218,g4267,I5720,g2390,g2397,g5199,g1046,g2505,
    g3788,g6034,g6434,I6299,g4438,I5750,I2929,g6347,g1191,g3192,I3746,g5947,
    g3485,g1637,g2631,I8656,g3854,g6445,g2817,g4519,g6413,I8249,I5790,I6078,
    g4387,I6340,g5923,I3468,g1802,I6959,g3219,I4318,I7634,g5727,I5427,g3726,
    g3031,g6117,g5880,g1642,g6482,I5904,g3749,g5886,g6657,I3152,g1334,I2053,
    g5114,I5403,g5314,I6972,I2453,g1654,I5529,g3975,g3911,I5148,g6581,g1880,
    g1603,I5618,g2772,g2743,g6784,g2890,g1875,I4300,g1978,g1387,g3796,g1659,
    I3629,g3124,g2856,g2010,g2734,I3902,g4524,g836,g3540,g5887,g1542,g3177,
    I3717,I6895,I5542,g4577,g4717,g4465,g5433,g3742,g5017,g2863,g3199,g5550,
    g3781,g5891,g3898,g3900,g1118,g3797,g6850,g6163,g5726,g3510,g3910,I5457,
    g2688,g2857,g3291,g2976,I2402,I6923,g1056,g3502,g1529,g3984,g1649,g1348,
    g5248,g4636,I2394,g5255,I9031,g2760,g3488,g6709,I4587,I6733,I7487,g4187,
    I5591,I9005,g3886,g2779,g4904,g4812,g1279,g1111,g5112,g2588,g6449,I6769,
    g4763,g3136,g2739,g1549,g947,g6894,I9149,I5851,g3739,g4536,g6735,I2970,
    g858,I3115,I3251,g6303,g3465,g3322,g3783,g4522,g6440,g2043,I3158,g6039,
    I8764,g3096,I4343,g3851,g1552,I8617,g850,g5576,g4537,g4410,g5149,g6276,
    g4612,g2914,g6616,I2376,g3342,g4328,g4092,g4351,I7963,g3481,g2820,g2936,
    g2026,g3354,I5204,g5119,g5701,g1358,g5577,g4213,g6120,g2922,I6812,g6788,
    g5893,g2908,g6095,g2060,g6617,g6906,g5975,g5821,g4512,g6702,g3001,g4166,
    g6516,g6409,I3148,g3761,g4529,g4773,g3830,g2079,g4155,g6892,g6936,I2955,
    g2840,g3745,g5544,g4450,g1559,I6069,g4463,g943,I8837,g6078,g5061,I6701,
    g6478,g866,g6035,g4720,g3677,g3140,g2954,g2966,g5046,g6656,g4193,g2032,
    g1749,g3814,g5391,g2568,g2912,g5467,g2357,g1323,g4625,g4232,g1666,g4938,
    g5019,g6236,g6295,g5684,g1528,g1351,g5115,g5251,g5069,g5315,I5094,g1655,
    g1410,g5167,g6899,g929,g5385,g2778,g3370,g2894,I7007,g4163,g4525,g3483,
    g6194,g1829,g5542,g3306,g2998,g4158,g1555,g3790,g2039,g3187,g3387,g3461,
    g4587,I6033,g4179,g5554,g5455,g3904,g3200,g2919,g2952,g4455,g3599,g4545,
    g4416,g5090,g4020,g6212,I7910,g5456,g5649,g4507,g2764,g6430,g5155,g3016,
    g6229,g5260,g6289,g4628,g4515,g2120,g6479,g2906,g2789,g5118,g2771,g6620,
    g5193,g4967,I5360,g3532,g3536,g3539,g3544,g5598,g6249,g4666,g4630,g4627,
    g3629,g3328,g6085,g4648,g4407,g5232,g2340,g5938,g5909,g3554,g2941,g3903,
    g1474,g6640,g6549,g4172,g3930,g4372,g3490,g4667,g4653,g4651,g3166,g3366,
    g6829,g3649,g6911,g3155,g3698,g6270,g4792,g1417,g4471,g6473,g6397,g1628,
    g4621,g3953,g5158,g4993,g6124,g6324,g3880,g2121,g6394,g3279,g3619,g3167,
    g5311,g5013,g4468,g3367,g3652,g3843,g3533,g4593,g4277,g3686,g5180,g4950,
    g5380,g4160,g3923,g3321,g2089,g6245,g3670,g3625,I5359,g5559,g5024,g6144,
    g6344,g6272,g2948,g2137,g6259,g2955,g6088,g6852,g6847,g6923,g6918,g6917,
    g5515,g5364,g1499,g4835,g3687,g4271,g4004,g4611,g3985,g4300,g3341,g6650,
    g4541,g4199,g3645,g5123,g4670,g3691,g4209,g3816,g4353,g3989,g6336,g6246,
    g6768,g6750,g4744,g3434,g3659,g5351,g5326,g3358,g5648,g6934,g3275,g3311,
    g5410,g3615,g2062,g3374,g4600,g4054,g6096,g1436,g5172,g4877,g3180,g5618,
    g5506,g5143,g6913,g5235,g4580,g2085,g6266,g5555,g5014,g2166,g6248,g6342,
    g6264,g5621,g5508,g3628,g6255,g6081,g3630,g6692,g3300,g6154,g6354,g4184,
    g3934,g5494,g5443,g4384,g4339,g3971,g4838,g3123,g3323,g4672,g4635,g4631,
    g2733,g3666,g6129,g6329,g3888,g2073,g5360,g6828,g4285,g3351,g6830,g3648,
    g3655,g1706,g6068,g4044,g6468,g1609,g3172,g3278,g3372,g2781,g3618,g3667,
    g3143,g3282,g6716,g6682,g6149,g3693,g3134,g3334,g6848,g3741,g6843,g5153,
    g5209,g5353,g5327,g6241,g1808,g3113,g5558,g5018,g6644,g6152,g6258,g4178,
    g3959,g1575,g4378,g4831,g5492,g5441,g5600,g5502,g6614,g6556,g4947,g3360,
    g6125,g1419,g918,g3641,g4873,g4037,g2896,g4495,g3913,g3379,g5175,g5094,
    g3658,g6061,g5500,g5430,g5074,g3611,g4042,g5184,g4442,g4239,g4164,g3958,
    g2807,g5424,g6145,g3997,g3425,g3694,g6345,g6273,g3132,g3680,g6637,g3353,
    g2142,g2255,g6159,g2081,g3558,g5499,g5451,g4389,g4171,g3956,g6315,g3849,
    g4371,g4429,g4253,g4787,g2937,g6047,g6874,g6873,g2267,g1716,g5444,g1574,
    g5269,g4684,g4584,g4791,g3936,g6243,g6935,g2746,g4759,g4500,g6128,g5414,
    g6130,g5660,g3375,g4449,g4266,g3651,g4865,g4776,g2953,g2068,g3285,g4833,
    g5178,g5679,g5378,g3339,g1689,g5182,g2699,g2747,g6090,g4362,g3996,g3672,
    g4052,g3643,g4452,g3820,g6056,g1826,g6148,g6348,g5560,g5044,g3634,g6155,
    g6851,g6846,g3551,g3099,g3304,g4486,g3499,g4730,g5632,g5095,g4794,g6260,
    g5495,g1138,g3613,g6318,g3865,g901,g5164,g5194,g5233,g2821,g5454,g4549,
    g5553,g5012,g6321,g3873,g3660,g6625,g4045,g4445,g4235,g6253,g4373,g4001,
    g5189,g4491,g6909,g4169,g3966,g5171,g4369,g3999,g3679,g4602,g5371,g3378,
    g5429,g5956,g5783,g4868,g4774,g5675,g3135,g4459,g4245,g3335,g3831,g3182,
    g3288,g3382,g4793,g4015,g2107,g6141,g6341,g6261,g6645,g3632,g3437,g2853,
    g3653,g5201,g4859,g3208,g2551,g3302,g6158,g5449,g5246,g5604,g5098,g4021,
    g5498,g1585,g6275,g6311,g3837,g4671,g4645,g4641,g4247,g4007,g4826,g5162,
    g5088,g5362,g3296,g5419,g2935,g6559,g5728,g5623,g5486,g5185,g3171,g3371,
    g6628,g2138,g4165,g3927,g4048,g4448,g3815,g3281,g4827,g4333,g3964,I2566,
    g1633,g3684,g4396,g3338,g2056,g5406,g3309,g5635,g5682,g5487,g6123,g6323,
    g3877,g3759,g5226,g6151,g3449,g6648,g5173,g5373,g4181,g3939,g2720,g4685,
    g4591,g5169,g5093,g5369,I4040,g3362,g6343,g6268,g6693,g6334,g3858,g6555,
    g2909,g2092,g4041,g6313,g3841,g5940,g4673,g4656,g4654,g5188,g6908,g6907,
    g5216,g6094,g4168,g3925,g4368,g3998,g5671,g3678,g5428,g4058,g3635,g2860,
    g3682,g3305,g2960,g5910,g5816,g3755,g2659,g1686,g5883,g3373,g5217,g4866,
    g4863,g4777,g3283,g3602,I2574,g5165,g6777,g6762,g3718,g1157,g3767,g4688,
    g4568,g1784,g2021,g6799,g4948,g6782,g2794,g3203,g6132,g6238,g6153,g4183,
    g3965,g4383,g6558,g5181,g3689,g4588,g2419,g5197,g4161,g3931,g4361,g3995,
    g3671,g4051,g6092,g2323,g5562,g5228,g3609,g6262,g6736,g3758,g4043,g3365,
    g1558,g5673,g4347,g3986,g3133,g3333,g3774,g4697,g4589,g3780,g6737,g6077,
    g3662,g6643,g3290,g6634,g6545,g2113,g1576,g6099,g3181,g3381,g3685,g3700,
    g3421,g2846,g5569,g5348,g4597,g6613,g6554,g4739,g2850,g6269,g4937,g4668,
    g4642,g4638,g3631,g2160,g4390,g3301,g4156,g3926,g4942,g5183,g5023,g3935,
    g4363,g4032,g4053,g4453,g4238,g5161,g3669,g5361,g3368,g6135,g5665,g6831,
    g4544,g6288,g4357,g3990,g5146,g6916,g5633,g6749,g6798,g4946,g6781,g5944,
    g5778,g5240,g5043,g3941,g2307,g6302,g6719,g1570,g4683,g4585,g5681,g3688,
    g4735,g2018,g6265,g4782,g4661,g4637,g4634,g4949,g3326,g6770,g6754,g3760,
    g5936,g4039,g5317,g3383,g5601,g3608,g3924,g4583,g3161,g2339,g3361,g4616,
    g4231,g3665,g3127,g3327,g3146,g3633,g5937,g5775,g3103,g3303,g5668,g6338,
    g6251,g5190,g5501,g5156,g5356,g5265,g5942,g4789,g3316,g5954,g5163,g6098,
    g3147,g5363,g3681,g5053,g4599,g3697,g5157,g5357,g4244,g4340,g3972,g3117,
    g3317,g4035,g6086,g4214,g1822,g1620,g3784,g2916,g3479,g6131,g3668,g6331,
    g3891,g4236,g3907,g3294,g5949,g3190,g6766,g3156,g3356,g5646,g2873,g1845,
    g6748,g5603,g5504,g5484,g4928,g3704,g4464,g4272,g4785,g6091,g3810,g5952,
    g5616,g5505,g6718,g6767,g3157,g3357,g4489,g2770,g5503,g3626,g4038,g5617,
    g3683,g4836,g3661,g6247,g3627,g5945,g2808,g2009,g3292,g3646,g2759,g6910,
    g3603,g3484,g5482,g3702,g6066,g5214,g3616,g6055,g6133,g5663,g6333,g3896,
    g3764,g5402,g5236,g4708,g5556,g5015,g3277,g3617,g6093,g2897,g6256,g6816,
    g4829,g6263,g4874,g3709,g5557,g5016,g3340,g6631,g3522,g4177,g3933,g5948,
    g5779,g4377,g3690,g5955,g5782,g5350,g5325,g5438,g5224,g2868,g1316,g3310,
    g4797,g5212,g3663,g2793,g2015,g4344,g3981,g5229,g6772,g3762,g4694,g1481,
    g4578,g3657,g2721,g4488,g4701,g4596,g3928,g3899,g3464,g5620,g5507,g4870,
    g4779,g3295,g2671,g2263,g3089,g3489,g2607,g5192,g5485,g5941,g5777,g4230,
    g3756,g6126,g6326,g3833,g4033,g2758,g3350,g6924,g6920,g6919,g5176,g4395,
    g5376,g5911,g5817,g6127,g6327,g3884,g5225,g4342,g3978,g6146,g6346,g6274,
    g4354,I5352,g3529,g3531,g3535,g3538,g5177,g6240,g4205,g3620,g1027,g2685,
    g2700,g6316,g3855,g5898,g5800,g4401,g1514,g5900,g5804,g2950,g2156,g5245,
    g1763,g4828,g3298,g4830,g5144,g4592,g6914,g2101,g5488,g4932,g1416,g5683,
    g6317,g3862,g5215,g4864,g5951,g5780,g4677,g4652,g4646,g3176,g3376,g3286,
    g3765,g4349,g6060,g3518,g3521,g3526,g3530,g3610,g6739,g3324,g6079,g5122,
    g3377,g4352,g3988,g4867,g4811,g6156,g3287,g5096,g4186,g3973,g5496,g5446,
    g6250,g4280,g3144,g3344,g5142,g3819,g6912,g6157,g5481,g3701,g5497,g5447,
    g5154,g5354,g5249,g4461,g4241,g4756,I5351,g5218,g3650,g4345,g3982,g3336,
    g4359,g3806,g2024,g3905,g3887,g3276,g3122,g2435,g2732,g4047,g6646,g3433,
    g905,g5953,g5781,g6084,g6603,g5677,g3195,g3337,g5349,g5324,g5198,g5398,
    g6647,g1691,g3692,g3154,g4800,g5152,g6320,g3869,g5211,g4860,g5186,g5599,
    g4490,g3293,g6771,g6758,g3329,g5170,g5091,g4456,g3829,g4348,g3987,g4355,
    g5939,g5776,g2294,g4698,g4586,g5483,g3703,g6738,g6244,g2356,g6140,g6340,
    g6257,g5187,g6082,g4057,g5904,g5812,g5200,g4457,g4261,g5241,g3349,g2053,
    g5145,g6915,g4834,g4686,g4590,g5191,g3699,g4598,g5637,g5159,g5359,g3644,
    g3319,g3352,g5047,g3954,g2311,g3186,g3170,g3614,g3325,g4341,g3977,g2782,
    g3280,g4691,g4581,g5935,g2949,g3511,g3517,g3520,g3525,g5234,g3636,g2292,
    g6089,g6731,g6717,g4427,g6557,g4358,g3991,g2084,g5213,g4862,g6254,g6150,
    g5902,g5808,g3145,g3345,g6773,g3763,g3191,g4180,g3929,g5166,g3637,g4832,
    g6769,g3307,g3359,g3757,g3315,g3642,g3654,g5619,I8376,I8393,I8394,I8395,
    I8377,g5659,g2100,g1582,g5374,g3598,I8136,g5666,I8137,g6280,I9057,I8081,
    I9064,I9065,I9066,g5372,I8129,I8367,I8368,I8369,I8370,g4243,g5202,g4000,
    I8349,I8345,I8346,I8347,I8348,g6703,I8119,g5674,g6747,I8211,I8386,g5680,
    g6358,I8387,g6281,I8385,I8359,g4233,g5672,g5048,I8128,I7970,I7987,I8118,
    g1589,I8358,g6659,g6073,g6741,g6929,g3992,g5678,g2080,I7980,I8360,I8356,
    I8357,I8379,g6357,g5066,I8209,g5662,I7972,I9059,g6279,g5669,g5368,I7979,
    g4936,g6926,I8378,I8135,g3012,g6400,g6927,g6660,I8208,g3028,I8138,I9058,
    g5060,g4819,I7978,I7989,I7971,g3215,I8774,g3503,I7969,g4941,I7988,I8080,
    g6669,I8126,g5062,g6359,I8779,I7981,I8127,I8778,I8210,g5377,I8117,I8079,
    g6335,g5065,g2995,g2095,g1573,g6683,g5676,I8773,g4432,g5068,I7990,I8120,
    g2067,g4234,g5227,I8082,g5370,g3013,g6740,g6928,g2951,g6705,g6075,g5367,
    I7217,I7216,I7571,I7569,I2073,I2072,I2796,I2795,g948,I2014,I2015,I4205,
    I4203,I3875,I3874,g3109,I5536,I5537,I5658,g3983,I5657,I2527,I2528,I4444,
    I5271,I5269,I2898,I2897,I2797,I2245,I2244,I3988,I2543,I2544,I1963,I1961,
    I5209,I5207,I7562,I7231,I7232,I6744,I6745,I4182,I6186,g4301,I6185,I7441,
    I7439,I6026,g4223,g4221,I2768,I2766,I3933,g2731,I3894,I3895,I7238,I7239,
    I4160,I4161,I2934,I2933,I3179,I3177,I6187,g3955,I6027,I4233,g2769,I3953,
    I3954,g1044,I2081,I2082,g4674,I6391,g4504,I6390,g4680,I2080,I8195,I8194,
    g1534,I2498,I2499,I2497,g1042,g1036,g939,I1987,I1988,I2061,I2062,I2676,
    I2674,I2767,I7528,I7529,I7434,I7432,I2074,I7210,I7208,I6964,I6962,I5208,
    I5302,I5300,I7535,I7536,I6195,I6196,I2542,I1994,I4445,I2060,I5189,I5187,
    I3178,I4920,I4919,I2003,I3916,I3914,I5309,I5307,I5759,I6659,g4762,I4940,
    I4939,I2935,I3412,I3413,I3411,I3189,I3188,I3990,I4151,I4152,I2090,I2089,
    g5862,I9050,I5766,g3961,g3957,g3968,I5227,I5228,I7527,I5226,g4049,I7224,
    I7223,I5767,I5535,g2944,I4921,I6028,I7244,I5188,I5270,I9051,I9052,I5308,
    I2506,g1047,I3445,I3169,I3170,g1540,I3168,I7556,I7555,I5196,I5195,I7563,
    I7440,I2507,I1995,I3446,I3447,I7237,g2757,I3934,I3935,I6743,I4183,I7557,
    I2300,I2299,I5197,I4159,I3741,I3739,I6660,I6661,I5257,I2526,I5301,I4204,
    I7218,I6175,I3455,I6500,I6499,I3846,I4210,I6474,I6475,g2698,I3847,I3848,
    g1518,I7520,I4784,I4782,I1952,I1951,I8202,I8201,I1986,I5760,I5768,I1970,
    I1969,I7225,I7209,I2301,I7245,I3740,I6963,I3456,I3457,I3126,I3125,I3400,
    I3398,I4526,I4527,I4528,g2795,I6176,I6177,I7230,I7433,I3127,I4234,I4235,
    I5784,I5782,I7550,I7548,I4546,I4545,I5294,I5292,g937,I1979,I1980,g4472,
    g1473,g1470,g1459,g928,I1962,I7097,I4547,I3697,I7312,I7311,I2109,I2110,
    I2013,g2804,I4009,I4010,g5863,I2022,I2021,I7576,g5688,I3190,I3952,I7549,
    I7577,I5647,g3974,I1978,I7246,I4150,g3621,I4008,I2675,g926,I1953,I3893,
    I4212,I7313,I2108,I5244,I5242,I7534,I7522,I7521,I6194,I3970,I4941,g3979,
    I7542,I7541,I2682,I2681,I4211,I3876,I2091,I3915,I4783,I7543,g930,I1971,
    I7570,I5293,I2246,I6392,g944,I2004,I2005,I6473,g2719,I8203,I2899,g941,
    I1996,I2508,g2745,g2791,I3989,I8196,I5259,g1560,g4610,I6501,I3399,I3698,
    I3699,g950,I2023,I4446,I5783,g2940,I5761,I3972,I7098,I7099,g2780,I3971,
    I5258,I7564,I5648,I5649,I5243,I2683,I7578,I5659,I4184,g3528,g3664,g3656,
    g3647,g1449,g1418,g1879;

  //scan intermediate wires
  wire tdo_0  ;
  wire tdo_1  ;
  wire tdo_2  ;
  wire tdo_3  ;
  wire tdo_4  ;
  wire tdo_5  ;
  wire tdo_6  ;
  wire tdo_7  ;
  wire tdo_8  ;
  wire tdo_9  ;
  wire tdo_10 ;
  wire tdo_11 ;
  wire tdo_12 ;
  wire tdo_13 ;
  wire tdo_14 ;
  wire tdo_15 ;
  wire tdo_16 ;
  wire tdo_17 ;
  wire tdo_18 ;
  wire tdo_19 ;
  wire tdo_20 ;
  wire tdo_21 ;
  wire tdo_22 ;
  wire tdo_23 ;
  wire tdo_24 ;
  wire tdo_25 ;
  wire tdo_26 ;
  wire tdo_27 ;
  wire tdo_28 ;
  wire tdo_29 ;
  wire tdo_30 ;
  wire tdo_31 ;
  wire tdo_32 ;
  wire tdo_33 ;
  wire tdo_34 ;
  wire tdo_35 ;
  wire tdo_36 ;
  wire tdo_37 ;
  wire tdo_38 ;
  wire tdo_39 ;
  wire tdo_40 ;
  wire tdo_41 ;
  wire tdo_42 ;
  wire tdo_43 ;
  wire tdo_44 ;
  wire tdo_45 ;
  wire tdo_46 ;
  wire tdo_47 ;
  wire tdo_48 ;
  wire tdo_49 ;
  wire tdo_50 ;
  wire tdo_51 ;
  wire tdo_52 ;
  wire tdo_53 ;
  wire tdo_54 ;
  wire tdo_55 ;
  wire tdo_56 ;
  wire tdo_57 ;
  wire tdo_58 ;
  wire tdo_59 ;
  wire tdo_60 ;
  wire tdo_61 ;
  wire tdo_62 ;
  wire tdo_63 ;
  wire tdo_64 ;
  wire tdo_65 ;
  wire tdo_66 ;
  wire tdo_67 ;
  wire tdo_68 ;
  wire tdo_69 ;
  wire tdo_70 ;
  wire tdo_71 ;
  wire tdo_72 ;
  wire tdo_73 ;
  wire tdo_74 ;
  wire tdo_75 ;
  wire tdo_76 ;
  wire tdo_77 ;
  wire tdo_78 ;
  wire tdo_79 ;
  wire tdo_80 ;
  wire tdo_81 ;
  wire tdo_82 ;
  wire tdo_83 ;
  wire tdo_84 ;
  wire tdo_85 ;
  wire tdo_86 ;
  wire tdo_87 ;
  wire tdo_88 ;
  wire tdo_89 ;
  wire tdo_90 ;
  wire tdo_91 ;
  wire tdo_92 ;
  wire tdo_93 ;
  wire tdo_94 ;
  wire tdo_95 ;
  wire tdo_96 ;
  wire tdo_97 ;
  wire tdo_98 ;
  wire tdo_99 ;
  wire tdo_100;
  wire tdo_101;
  wire tdo_102;
  wire tdo_103;
  wire tdo_104;
  wire tdo_105;
  wire tdo_106;
  wire tdo_107;
  wire tdo_108;
  wire tdo_109;
  wire tdo_110;
  wire tdo_111;
  wire tdo_112;
  wire tdo_113;
  wire tdo_114;
  wire tdo_115;
  wire tdo_116;
  wire tdo_117;
  wire tdo_118;
  wire tdo_119;
  wire tdo_120;
  wire tdo_121;
  wire tdo_122;
  wire tdo_123;
  wire tdo_124;
  wire tdo_125;
  wire tdo_126;
  wire tdo_127;
  wire tdo_128;
  wire tdo_129;
  wire tdo_130;
  wire tdo_131;
  wire tdo_132;
  wire tdo_133;
  wire tdo_134;
  wire tdo_135;
  wire tdo_136;
  wire tdo_137;
  wire tdo_138;
  wire tdo_139;
  wire tdo_140;
  wire tdo_141;
  wire tdo_142;
  wire tdo_143;
  wire tdo_144;
  wire tdo_145;
  wire tdo_146;
  wire tdo_147;
  wire tdo_148;
  wire tdo_149;
  wire tdo_150;
  wire tdo_151;
  wire tdo_152;
  wire tdo_153;
  wire tdo_154;
  wire tdo_155;
  wire tdo_156;
  wire tdo_157;
  wire tdo_158;
  wire tdo_159;
  wire tdo_160;
  wire tdo_161;
  wire tdo_162;
  wire tdo_163;
  wire tdo_164;
  wire tdo_165;
  wire tdo_166;
  wire tdo_167;
  wire tdo_168;
  wire tdo_169;
  wire tdo_170;
  wire tdo_171;
  wire tdo_172;
  wire tdo_173;
  wire tdo_174;
  wire tdo_175;
  wire tdo_176;
  wire tdo_177;
  wire tdo_178;
  wire tdo_179;
  wire tdo_180;
  wire tdo_181;
  wire tdo_182;
  wire tdo_183;
  wire tdo_184;
  wire tdo_185;
  wire tdo_186;
  wire tdo_187;
  wire tdo_188;
  wire tdo_189;
  wire tdo_190;
  wire tdo_191;
  wire tdo_192;
  wire tdo_193;
  wire tdo_194;
  wire tdo_195;
  wire tdo_196;
  wire tdo_197;
  wire tdo_198;
  wire tdo_199;
  wire tdo_200;
  wire tdo_201;
  wire tdo_202;
  wire tdo_203;
  wire tdo_204;
  wire tdo_205;
  wire tdo_206;
  wire tdo_207;
  wire tdo_208;
  wire tdo_209;

  int_SFF_XXXX SFF_0   (bistsel,TDO_ISR,TDI_ISR,int_hold,g4130,CK,clockdr,updatedr,shiftdr,tdo_0  ,g678);
  int_SFF_XXXX SFF_1   (bistsel,TDO_ISR,tdo_0  ,int_hold,g6823,CK,clockdr,updatedr,shiftdr,tdo_1  ,g332);
  int_SFF_XXXX SFF_2   (bistsel,TDO_ISR,tdo_1  ,int_hold,g6940,CK,clockdr,updatedr,shiftdr,tdo_2  ,g123);
  int_SFF_XXXX SFF_3   (bistsel,TDO_ISR,tdo_2  ,int_hold,g6102,CK,clockdr,updatedr,shiftdr,tdo_3  ,g207);
  int_SFF_XXXX SFF_4   (bistsel,TDO_ISR,tdo_3  ,int_hold,g4147,CK,clockdr,updatedr,shiftdr,tdo_4  ,g695);
  int_SFF_XXXX SFF_5   (bistsel,TDO_ISR,tdo_4  ,int_hold,g4841,CK,clockdr,updatedr,shiftdr,tdo_5  ,g461);
  int_SFF_XXXX SFF_6   (bistsel,TDO_ISR,tdo_5  ,int_hold,g6725,CK,clockdr,updatedr,shiftdr,tdo_6  ,g18);
  int_SFF_XXXX SFF_7   (bistsel,TDO_ISR,tdo_6  ,int_hold,g3232,CK,clockdr,updatedr,shiftdr,tdo_7  ,g292);
  int_SFF_XXXX SFF_8   (bistsel,TDO_ISR,tdo_7  ,int_hold,g4119,CK,clockdr,updatedr,shiftdr,tdo_8  ,g331);
  int_SFF_XXXX SFF_9   (bistsel,TDO_ISR,tdo_8  ,int_hold,g4141,CK,clockdr,updatedr,shiftdr,tdo_9  ,g689);
  int_SFF_XXXX SFF_10  (bistsel,TDO_ISR,tdo_9  ,int_hold,g6726,CK,clockdr,updatedr,shiftdr,tdo_10 ,g24);
  int_SFF_XXXX SFF_11  (bistsel,TDO_ISR,tdo_10 ,int_hold,g6507,CK,clockdr,updatedr,shiftdr,tdo_11 ,g465);
  int_SFF_XXXX SFF_12  (bistsel,TDO_ISR,tdo_11 ,int_hold,g6590,CK,clockdr,updatedr,shiftdr,tdo_12 ,g84);
  int_SFF_XXXX SFF_13  (bistsel,TDO_ISR,tdo_12 ,int_hold,g3231,CK,clockdr,updatedr,shiftdr,tdo_13 ,g291);
  int_SFF_XXXX SFF_14  (bistsel,TDO_ISR,tdo_13 ,int_hold,g5330,CK,clockdr,updatedr,shiftdr,tdo_14 ,g676);
  int_SFF_XXXX SFF_15  (bistsel,TDO_ISR,tdo_14 ,int_hold,g5147,CK,clockdr,updatedr,shiftdr,tdo_15 ,g622);
  int_SFF_XXXX SFF_16  (bistsel,TDO_ISR,tdo_15 ,int_hold,g4839,CK,clockdr,updatedr,shiftdr,tdo_16 ,g117);
  int_SFF_XXXX SFF_17  (bistsel,TDO_ISR,tdo_16 ,int_hold,g6105,CK,clockdr,updatedr,shiftdr,tdo_17 ,g278);
  int_SFF_XXXX SFF_18  (bistsel,TDO_ISR,tdo_17 ,int_hold,g5138,CK,clockdr,updatedr,shiftdr,tdo_18 ,g128);
  int_SFF_XXXX SFF_19  (bistsel,TDO_ISR,tdo_18 ,int_hold,g4122,CK,clockdr,updatedr,shiftdr,tdo_19 ,g598);
  int_SFF_XXXX SFF_20  (bistsel,TDO_ISR,tdo_19 ,int_hold,g6827,CK,clockdr,updatedr,shiftdr,tdo_20 ,g554);
  int_SFF_XXXX SFF_21  (bistsel,TDO_ISR,tdo_20 ,int_hold,g6745,CK,clockdr,updatedr,shiftdr,tdo_21 ,g496);
  int_SFF_XXXX SFF_22  (bistsel,TDO_ISR,tdo_21 ,int_hold,g6405,CK,clockdr,updatedr,shiftdr,tdo_22 ,g179);
  int_SFF_XXXX SFF_23  (bistsel,TDO_ISR,tdo_22 ,int_hold,g6729,CK,clockdr,updatedr,shiftdr,tdo_23 ,g48);
  int_SFF_XXXX SFF_24  (bistsel,TDO_ISR,tdo_23 ,int_hold,g6595,CK,clockdr,updatedr,shiftdr,tdo_24 ,g590);
  int_SFF_XXXX SFF_25  (bistsel,TDO_ISR,tdo_24 ,int_hold,g6826,CK,clockdr,updatedr,shiftdr,tdo_25 ,g551);
  int_SFF_XXXX SFF_26  (bistsel,TDO_ISR,tdo_25 ,int_hold,g4134,CK,clockdr,updatedr,shiftdr,tdo_26 ,g682);
  int_SFF_XXXX SFF_27  (bistsel,TDO_ISR,tdo_26 ,int_hold,g6599,CK,clockdr,updatedr,shiftdr,tdo_27 ,g11);
  int_SFF_XXXX SFF_28  (bistsel,TDO_ISR,tdo_27 ,int_hold,g4857,CK,clockdr,updatedr,shiftdr,tdo_28 ,g606);
  int_SFF_XXXX SFF_29  (bistsel,TDO_ISR,tdo_28 ,int_hold,g6406,CK,clockdr,updatedr,shiftdr,tdo_29 ,g188);
  int_SFF_XXXX SFF_30  (bistsel,TDO_ISR,tdo_29 ,int_hold,g5148,CK,clockdr,updatedr,shiftdr,tdo_30 ,g646);
  int_SFF_XXXX SFF_31  (bistsel,TDO_ISR,tdo_30 ,int_hold,g4117,CK,clockdr,updatedr,shiftdr,tdo_31 ,g327);
  int_SFF_XXXX SFF_32  (bistsel,TDO_ISR,tdo_31 ,int_hold,g6582,CK,clockdr,updatedr,shiftdr,tdo_32 ,g361);
  int_SFF_XXXX SFF_33  (bistsel,TDO_ISR,tdo_32 ,int_hold,g3229,CK,clockdr,updatedr,shiftdr,tdo_33 ,g289);
  int_SFF_XXXX SFF_34  (bistsel,TDO_ISR,tdo_33 ,int_hold,g5700,CK,clockdr,updatedr,shiftdr,tdo_34 ,g398);
  int_SFF_XXXX SFF_35  (bistsel,TDO_ISR,tdo_34 ,int_hold,g4136,CK,clockdr,updatedr,shiftdr,tdo_35 ,g684);
  int_SFF_XXXX SFF_36  (bistsel,TDO_ISR,tdo_35 ,int_hold,g4858,CK,clockdr,updatedr,shiftdr,tdo_36 ,g619);
  int_SFF_XXXX SFF_37  (bistsel,TDO_ISR,tdo_36 ,int_hold,g5876,CK,clockdr,updatedr,shiftdr,tdo_37 ,g208);
  int_SFF_XXXX SFF_38  (bistsel,TDO_ISR,tdo_37 ,int_hold,g3239,CK,clockdr,updatedr,shiftdr,tdo_38 ,g248);
  int_SFF_XXXX SFF_39  (bistsel,TDO_ISR,tdo_38 ,int_hold,g5698,CK,clockdr,updatedr,shiftdr,tdo_39 ,g390);
  int_SFF_XXXX SFF_40  (bistsel,TDO_ISR,tdo_39 ,int_hold,g5328,CK,clockdr,updatedr,shiftdr,tdo_40 ,g625);
  int_SFF_XXXX SFF_41  (bistsel,TDO_ISR,tdo_40 ,int_hold,g4133,CK,clockdr,updatedr,shiftdr,tdo_41 ,g681);
  int_SFF_XXXX SFF_42  (bistsel,TDO_ISR,tdo_41 ,int_hold,g4847,CK,clockdr,updatedr,shiftdr,tdo_42 ,g437);
  int_SFF_XXXX SFF_43  (bistsel,TDO_ISR,tdo_42 ,int_hold,g5877,CK,clockdr,updatedr,shiftdr,tdo_43 ,g276);
  int_SFF_XXXX SFF_44  (bistsel,TDO_ISR,tdo_43 ,int_hold,g6597,CK,clockdr,updatedr,shiftdr,tdo_44 ,g3);
  int_SFF_XXXX SFF_45  (bistsel,TDO_ISR,tdo_44 ,int_hold,g4120,CK,clockdr,updatedr,shiftdr,tdo_45 ,g323);
  int_SFF_XXXX SFF_46  (bistsel,TDO_ISR,tdo_45 ,int_hold,g3235,CK,clockdr,updatedr,shiftdr,tdo_46 ,g224);
  int_SFF_XXXX SFF_47  (bistsel,TDO_ISR,tdo_46 ,int_hold,g4137,CK,clockdr,updatedr,shiftdr,tdo_47 ,g685);
  int_SFF_XXXX SFF_48  (bistsel,TDO_ISR,tdo_47 ,int_hold,g6407,CK,clockdr,updatedr,shiftdr,tdo_48 ,g43);
  int_SFF_XXXX SFF_49  (bistsel,TDO_ISR,tdo_48 ,int_hold,g5470,CK,clockdr,updatedr,shiftdr,tdo_49 ,g157);
  int_SFF_XXXX SFF_50  (bistsel,TDO_ISR,tdo_49 ,int_hold,g6841,CK,clockdr,updatedr,shiftdr,tdo_50 ,g282);
  int_SFF_LSFR SFF_51  (bistsel,TDO_ISR,tdo_50 ,int_hold,g4149,CK,clockdr,updatedr,shiftdr,tdo_51 ,g697);
  int_SFF_XXXX SFF_52  (bistsel,TDO_ISR,tdo_51 ,int_hold,g6101,CK,clockdr,updatedr,shiftdr,tdo_52 ,g206);
  int_SFF_XXXX SFF_53  (bistsel,TDO_ISR,tdo_52 ,int_hold,g4844,CK,clockdr,updatedr,shiftdr,tdo_53 ,g449);
  int_SFF_XXXX SFF_54  (bistsel,TDO_ISR,tdo_53 ,int_hold,g4113,CK,clockdr,updatedr,shiftdr,tdo_54 ,g118);
  int_SFF_XXXX SFF_55  (bistsel,TDO_ISR,tdo_54 ,int_hold,g6504,CK,clockdr,updatedr,shiftdr,tdo_55 ,g528);
  int_SFF_XXXX SFF_56  (bistsel,TDO_ISR,tdo_55 ,int_hold,g3224,CK,clockdr,updatedr,shiftdr,tdo_56 ,g284);
  int_SFF_XXXX SFF_57  (bistsel,TDO_ISR,tdo_56 ,int_hold,g4855,CK,clockdr,updatedr,shiftdr,tdo_57 ,g426);
  int_SFF_XXXX SFF_58  (bistsel,TDO_ISR,tdo_57 ,int_hold,g4424,CK,clockdr,updatedr,shiftdr,tdo_58 ,g634);
  int_SFF_XXXX SFF_59  (bistsel,TDO_ISR,tdo_58 ,int_hold,g5582,CK,clockdr,updatedr,shiftdr,tdo_59 ,g669);
  int_SFF_XXXX SFF_60  (bistsel,TDO_ISR,tdo_59 ,int_hold,g6502,CK,clockdr,updatedr,shiftdr,tdo_60 ,g520);
  int_SFF_XXXX SFF_61  (bistsel,TDO_ISR,tdo_60 ,int_hold,g6107,CK,clockdr,updatedr,shiftdr,tdo_61 ,g281);
  int_SFF_XXXX SFF_62  (bistsel,TDO_ISR,tdo_61 ,int_hold,g5472,CK,clockdr,updatedr,shiftdr,tdo_62 ,g175);
  int_SFF_LSFR SFF_63  (bistsel,TDO_ISR,tdo_62 ,int_hold,g6602,CK,clockdr,updatedr,shiftdr,tdo_63 ,g15);
  int_SFF_XXXX SFF_64  (bistsel,TDO_ISR,tdo_63 ,int_hold,g5581,CK,clockdr,updatedr,shiftdr,tdo_64 ,g631);
  int_SFF_XXXX SFF_65  (bistsel,TDO_ISR,tdo_64 ,int_hold,g6587,CK,clockdr,updatedr,shiftdr,tdo_65 ,g69);
  int_SFF_XXXX SFF_66  (bistsel,TDO_ISR,tdo_65 ,int_hold,g4145,CK,clockdr,updatedr,shiftdr,tdo_66 ,g693);
  int_SFF_XXXX SFF_67  (bistsel,TDO_ISR,tdo_66 ,int_hold,g2585,CK,clockdr,updatedr,shiftdr,tdo_67 ,g337);
  int_SFF_XXXX SFF_68  (bistsel,TDO_ISR,tdo_67 ,int_hold,g4842,CK,clockdr,updatedr,shiftdr,tdo_68 ,g457);
  int_SFF_XXXX SFF_69  (bistsel,TDO_ISR,tdo_68 ,int_hold,g2586,CK,clockdr,updatedr,shiftdr,tdo_69 ,g486);
  int_SFF_XXXX SFF_70  (bistsel,TDO_ISR,tdo_69 ,int_hold,g1291,CK,clockdr,updatedr,shiftdr,tdo_70 ,g471);
  int_SFF_XXXX SFF_71  (bistsel,TDO_ISR,tdo_70 ,int_hold,g4118,CK,clockdr,updatedr,shiftdr,tdo_71 ,g328);
  int_SFF_XXXX SFF_72  (bistsel,TDO_ISR,tdo_71 ,int_hold,g3225,CK,clockdr,updatedr,shiftdr,tdo_72 ,g285);
  int_SFF_XXXX SFF_73  (bistsel,TDO_ISR,tdo_72 ,int_hold,g4853,CK,clockdr,updatedr,shiftdr,tdo_73 ,g418);
  int_SFF_XXXX SFF_74  (bistsel,TDO_ISR,tdo_73 ,int_hold,g4849,CK,clockdr,updatedr,shiftdr,tdo_74 ,g402);
  int_SFF_XXXX SFF_75  (bistsel,TDO_ISR,tdo_74 ,int_hold,g6512,CK,clockdr,updatedr,shiftdr,tdo_75 ,g297);
  int_SFF_XXXX SFF_76  (bistsel,TDO_ISR,tdo_75 ,int_hold,g3233,CK,clockdr,updatedr,shiftdr,tdo_76 ,g212);
  int_SFF_XXXX SFF_77  (bistsel,TDO_ISR,tdo_76 ,int_hold,g4851,CK,clockdr,updatedr,shiftdr,tdo_77 ,g410);
  int_SFF_XXXX SFF_78  (bistsel,TDO_ISR,tdo_77 ,int_hold,g4856,CK,clockdr,updatedr,shiftdr,tdo_78 ,g430);
  int_SFF_XXXX SFF_79  (bistsel,TDO_ISR,tdo_78 ,int_hold,g6854,CK,clockdr,updatedr,shiftdr,tdo_79 ,g33);
  int_SFF_XXXX SFF_80  (bistsel,TDO_ISR,tdo_79 ,int_hold,g1831,CK,clockdr,updatedr,shiftdr,tdo_80 ,g662);
  int_SFF_XXXX SFF_81  (bistsel,TDO_ISR,tdo_80 ,int_hold,g4843,CK,clockdr,updatedr,shiftdr,tdo_81 ,g453);
  int_SFF_XXXX SFF_82  (bistsel,TDO_ISR,tdo_81 ,int_hold,g6510,CK,clockdr,updatedr,shiftdr,tdo_82 ,g269);
  int_SFF_XXXX SFF_83  (bistsel,TDO_ISR,tdo_82 ,int_hold,g6591,CK,clockdr,updatedr,shiftdr,tdo_83 ,g574);
  int_SFF_XXXX SFF_84  (bistsel,TDO_ISR,tdo_83 ,int_hold,g4846,CK,clockdr,updatedr,shiftdr,tdo_84 ,g441);
  int_SFF_XXXX SFF_85  (bistsel,TDO_ISR,tdo_84 ,int_hold,g1288,CK,clockdr,updatedr,shiftdr,tdo_85 ,g664);
  int_SFF_XXXX SFF_86  (bistsel,TDO_ISR,tdo_85 ,int_hold,g5478,CK,clockdr,updatedr,shiftdr,tdo_86 ,g349);
  int_SFF_XXXX SFF_87  (bistsel,TDO_ISR,tdo_86 ,int_hold,g6840,CK,clockdr,updatedr,shiftdr,tdo_87 ,g211);
  int_SFF_XXXX SFF_88  (bistsel,TDO_ISR,tdo_87 ,int_hold,g6594,CK,clockdr,updatedr,shiftdr,tdo_88 ,g586);
  int_SFF_LSFR SFF_89  (bistsel,TDO_ISR,tdo_88 ,int_hold,g5580,CK,clockdr,updatedr,shiftdr,tdo_89 ,g571);
  int_SFF_XXXX SFF_90  (bistsel,TDO_ISR,tdo_89 ,int_hold,g6853,CK,clockdr,updatedr,shiftdr,tdo_90 ,g29);
  int_SFF_XXXX SFF_91  (bistsel,TDO_ISR,tdo_90 ,int_hold,g4840,CK,clockdr,updatedr,shiftdr,tdo_91 ,g326);
  int_SFF_XXXX SFF_92  (bistsel,TDO_ISR,tdo_91 ,int_hold,g4150,CK,clockdr,updatedr,shiftdr,tdo_92 ,g698);
  int_SFF_XXXX SFF_93  (bistsel,TDO_ISR,tdo_92 ,int_hold,g5490,CK,clockdr,updatedr,shiftdr,tdo_93 ,g654);
  int_SFF_XXXX SFF_94  (bistsel,TDO_ISR,tdo_93 ,int_hold,g6511,CK,clockdr,updatedr,shiftdr,tdo_94 ,g293);
  int_SFF_XXXX SFF_95  (bistsel,TDO_ISR,tdo_94 ,int_hold,g4142,CK,clockdr,updatedr,shiftdr,tdo_95 ,g690);
  int_SFF_XXXX SFF_96  (bistsel,TDO_ISR,tdo_95 ,int_hold,g4845,CK,clockdr,updatedr,shiftdr,tdo_96 ,g445);
  int_SFF_XXXX SFF_97  (bistsel,TDO_ISR,tdo_96 ,int_hold,g5694,CK,clockdr,updatedr,shiftdr,tdo_97 ,g374);
  int_SFF_XXXX SFF_98  (bistsel,TDO_ISR,tdo_97 ,int_hold,g6722,CK,clockdr,updatedr,shiftdr,tdo_98 ,g6);
  int_SFF_XXXX SFF_99  (bistsel,TDO_ISR,tdo_98 ,int_hold,g4139,CK,clockdr,updatedr,shiftdr,tdo_99 ,g687);
  int_SFF_XXXX SFF_100 (bistsel,TDO_ISR,tdo_99 ,int_hold,g5480,CK,clockdr,updatedr,shiftdr,tdo_100,g357);
  int_SFF_XXXX SFF_101 (bistsel,TDO_ISR,tdo_100,int_hold,g5697,CK,clockdr,updatedr,shiftdr,tdo_101,g386);
  int_SFF_XXXX SFF_102 (bistsel,TDO_ISR,tdo_101,int_hold,g6498,CK,clockdr,updatedr,shiftdr,tdo_102,g504);
  int_SFF_XXXX SFF_103 (bistsel,TDO_ISR,tdo_102,int_hold,g4126,CK,clockdr,updatedr,shiftdr,tdo_103,g665);
  int_SFF_XXXX SFF_104 (bistsel,TDO_ISR,tdo_103,int_hold,g5471,CK,clockdr,updatedr,shiftdr,tdo_104,g166);
  int_SFF_XXXX SFF_105 (bistsel,TDO_ISR,tdo_104,int_hold,g6505,CK,clockdr,updatedr,shiftdr,tdo_105,g541);
  int_SFF_XXXX SFF_106 (bistsel,TDO_ISR,tdo_105,int_hold,g6588,CK,clockdr,updatedr,shiftdr,tdo_106,g74);
  int_SFF_XXXX SFF_107 (bistsel,TDO_ISR,tdo_106,int_hold,g5475,CK,clockdr,updatedr,shiftdr,tdo_107,g338);
  int_SFF_XXXX SFF_108 (bistsel,TDO_ISR,tdo_107,int_hold,g4148,CK,clockdr,updatedr,shiftdr,tdo_108,g696);
  int_SFF_XXXX SFF_109 (bistsel,TDO_ISR,tdo_108,int_hold,g6501,CK,clockdr,updatedr,shiftdr,tdo_109,g516);
  int_SFF_XXXX SFF_110 (bistsel,TDO_ISR,tdo_109,int_hold,g6506,CK,clockdr,updatedr,shiftdr,tdo_110,g536);
  int_SFF_XXXX SFF_111 (bistsel,TDO_ISR,tdo_110,int_hold,g4135,CK,clockdr,updatedr,shiftdr,tdo_111,g683);
  int_SFF_XXXX SFF_112 (bistsel,TDO_ISR,tdo_111,int_hold,g5479,CK,clockdr,updatedr,shiftdr,tdo_112,g353);
  int_SFF_XXXX SFF_113 (bistsel,TDO_ISR,tdo_112,int_hold,g6824,CK,clockdr,updatedr,shiftdr,tdo_113,g545);
  int_SFF_LSFR SFF_114 (bistsel,TDO_ISR,tdo_113,int_hold,g3240,CK,clockdr,updatedr,shiftdr,tdo_114,g254);
  int_SFF_XXXX SFF_115 (bistsel,TDO_ISR,tdo_114,int_hold,g5476,CK,clockdr,updatedr,shiftdr,tdo_115,g341);
  int_SFF_XXXX SFF_116 (bistsel,TDO_ISR,tdo_115,int_hold,g3230,CK,clockdr,updatedr,shiftdr,tdo_116,g290);
  int_SFF_XXXX SFF_117 (bistsel,TDO_ISR,tdo_116,int_hold,g6721,CK,clockdr,updatedr,shiftdr,tdo_117,g2);
  int_SFF_XXXX SFF_118 (bistsel,TDO_ISR,tdo_117,int_hold,g3227,CK,clockdr,updatedr,shiftdr,tdo_118,g287);
  int_SFF_XXXX SFF_119 (bistsel,TDO_ISR,tdo_118,int_hold,g6925,CK,clockdr,updatedr,shiftdr,tdo_119,g336);
  int_SFF_XXXX SFF_120 (bistsel,TDO_ISR,tdo_119,int_hold,g5477,CK,clockdr,updatedr,shiftdr,tdo_120,g345);
  int_SFF_XXXX SFF_121 (bistsel,TDO_ISR,tdo_120,int_hold,g5489,CK,clockdr,updatedr,shiftdr,tdo_121,g628);
  int_SFF_XXXX SFF_122 (bistsel,TDO_ISR,tdo_121,int_hold,g4131,CK,clockdr,updatedr,shiftdr,tdo_122,g679);
  int_SFF_XXXX SFF_123 (bistsel,TDO_ISR,tdo_122,int_hold,g6727,CK,clockdr,updatedr,shiftdr,tdo_123,g28);
  int_SFF_XXXX SFF_124 (bistsel,TDO_ISR,tdo_123,int_hold,g4140,CK,clockdr,updatedr,shiftdr,tdo_124,g688);
  int_SFF_XXXX SFF_125 (bistsel,TDO_ISR,tdo_124,int_hold,g6842,CK,clockdr,updatedr,shiftdr,tdo_125,g283);
  int_SFF_XXXX SFF_126 (bistsel,TDO_ISR,tdo_125,int_hold,g4423,CK,clockdr,updatedr,shiftdr,tdo_126,g613);
  int_SFF_XXXX SFF_127 (bistsel,TDO_ISR,tdo_126,int_hold,g6723,CK,clockdr,updatedr,shiftdr,tdo_127,g10);
  int_SFF_XXXX SFF_128 (bistsel,TDO_ISR,tdo_127,int_hold,g6724,CK,clockdr,updatedr,shiftdr,tdo_128,g14);
  int_SFF_XXXX SFF_129 (bistsel,TDO_ISR,tdo_128,int_hold,g4132,CK,clockdr,updatedr,shiftdr,tdo_129,g680);
  int_SFF_XXXX SFF_130 (bistsel,TDO_ISR,tdo_129,int_hold,g6401,CK,clockdr,updatedr,shiftdr,tdo_130,g143);
  int_SFF_XXXX SFF_131 (bistsel,TDO_ISR,tdo_130,int_hold,g5491,CK,clockdr,updatedr,shiftdr,tdo_131,g672);
  int_SFF_XXXX SFF_132 (bistsel,TDO_ISR,tdo_131,int_hold,g4127,CK,clockdr,updatedr,shiftdr,tdo_132,g667);
  int_SFF_XXXX SFF_133 (bistsel,TDO_ISR,tdo_132,int_hold,g6278,CK,clockdr,updatedr,shiftdr,tdo_133,g366);
  int_SFF_XXXX SFF_134 (bistsel,TDO_ISR,tdo_133,int_hold,g6106,CK,clockdr,updatedr,shiftdr,tdo_134,g279);
  int_SFF_XXXX SFF_135 (bistsel,TDO_ISR,tdo_134,int_hold,g6744,CK,clockdr,updatedr,shiftdr,tdo_135,g492);
  int_SFF_LSFR SFF_136 (bistsel,TDO_ISR,tdo_135,int_hold,g6404,CK,clockdr,updatedr,shiftdr,tdo_136,g170);
  int_SFF_XXXX SFF_137 (bistsel,TDO_ISR,tdo_136,int_hold,g4138,CK,clockdr,updatedr,shiftdr,tdo_137,g686);
  int_SFF_XXXX SFF_138 (bistsel,TDO_ISR,tdo_137,int_hold,g3228,CK,clockdr,updatedr,shiftdr,tdo_138,g288);
  int_SFF_XXXX SFF_139 (bistsel,TDO_ISR,tdo_138,int_hold,g1289,CK,clockdr,updatedr,shiftdr,tdo_139,g638);
  int_SFF_XXXX SFF_140 (bistsel,TDO_ISR,tdo_139,int_hold,g4123,CK,clockdr,updatedr,shiftdr,tdo_140,g602);
  int_SFF_XXXX SFF_141 (bistsel,TDO_ISR,tdo_140,int_hold,g4658,CK,clockdr,updatedr,shiftdr,tdo_141,g642);
  int_SFF_XXXX SFF_142 (bistsel,TDO_ISR,tdo_141,int_hold,g5878,CK,clockdr,updatedr,shiftdr,tdo_142,g280);
  int_SFF_XXXX SFF_143 (bistsel,TDO_ISR,tdo_142,int_hold,g4125,CK,clockdr,updatedr,shiftdr,tdo_143,g663);
  int_SFF_XXXX SFF_144 (bistsel,TDO_ISR,tdo_143,int_hold,g4124,CK,clockdr,updatedr,shiftdr,tdo_144,g610);
  int_SFF_XXXX SFF_145 (bistsel,TDO_ISR,tdo_144,int_hold,g5874,CK,clockdr,updatedr,shiftdr,tdo_145,g148);
  int_SFF_XXXX SFF_146 (bistsel,TDO_ISR,tdo_145,int_hold,g6103,CK,clockdr,updatedr,shiftdr,tdo_146,g209);
  int_SFF_XXXX SFF_147 (bistsel,TDO_ISR,tdo_146,int_hold,g1294,CK,clockdr,updatedr,shiftdr,tdo_147,g675);
  int_SFF_XXXX SFF_148 (bistsel,TDO_ISR,tdo_147,int_hold,g1292,CK,clockdr,updatedr,shiftdr,tdo_148,g478);
  int_SFF_XXXX SFF_149 (bistsel,TDO_ISR,tdo_148,int_hold,g4115,CK,clockdr,updatedr,shiftdr,tdo_149,g122);
  int_SFF_XXXX SFF_150 (bistsel,TDO_ISR,tdo_149,int_hold,g6584,CK,clockdr,updatedr,shiftdr,tdo_150,g54);
  int_SFF_XXXX SFF_151 (bistsel,TDO_ISR,tdo_150,int_hold,g6596,CK,clockdr,updatedr,shiftdr,tdo_151,g594);
  int_SFF_XXXX SFF_152 (bistsel,TDO_ISR,tdo_151,int_hold,g3226,CK,clockdr,updatedr,shiftdr,tdo_152,g286);
  int_SFF_XXXX SFF_153 (bistsel,TDO_ISR,tdo_152,int_hold,g2587,CK,clockdr,updatedr,shiftdr,tdo_153,g489);
  int_SFF_XXXX SFF_154 (bistsel,TDO_ISR,tdo_153,int_hold,g4657,CK,clockdr,updatedr,shiftdr,tdo_154,g616);
  int_SFF_XXXX SFF_155 (bistsel,TDO_ISR,tdo_154,int_hold,g6589,CK,clockdr,updatedr,shiftdr,tdo_155,g79);
  int_SFF_XXXX SFF_156 (bistsel,TDO_ISR,tdo_155,int_hold,g3234,CK,clockdr,updatedr,shiftdr,tdo_156,g218);
  int_SFF_XXXX SFF_157 (bistsel,TDO_ISR,tdo_156,int_hold,g3238,CK,clockdr,updatedr,shiftdr,tdo_157,g242);
  int_SFF_XXXX SFF_158 (bistsel,TDO_ISR,tdo_157,int_hold,g6592,CK,clockdr,updatedr,shiftdr,tdo_158,g578);
  int_SFF_XXXX SFF_159 (bistsel,TDO_ISR,tdo_158,int_hold,g5473,CK,clockdr,updatedr,shiftdr,tdo_159,g184);
  int_SFF_XXXX SFF_160 (bistsel,TDO_ISR,tdo_159,int_hold,g4114,CK,clockdr,updatedr,shiftdr,tdo_160,g119);
  int_SFF_XXXX SFF_161 (bistsel,TDO_ISR,tdo_160,int_hold,g6800,CK,clockdr,updatedr,shiftdr,tdo_161,g668);
  int_SFF_XXXX SFF_162 (bistsel,TDO_ISR,tdo_161,int_hold,g5141,CK,clockdr,updatedr,shiftdr,tdo_162,g139);
  int_SFF_XXXX SFF_163 (bistsel,TDO_ISR,tdo_162,int_hold,g4854,CK,clockdr,updatedr,shiftdr,tdo_163,g422);
  int_SFF_XXXX SFF_164 (bistsel,TDO_ISR,tdo_163,int_hold,g6839,CK,clockdr,updatedr,shiftdr,tdo_164,g210);
  int_SFF_XXXX SFF_165 (bistsel,TDO_ISR,tdo_164,int_hold,g5699,CK,clockdr,updatedr,shiftdr,tdo_165,g394);
  int_SFF_XXXX SFF_166 (bistsel,TDO_ISR,tdo_165,int_hold,g3236,CK,clockdr,updatedr,shiftdr,tdo_166,g230);
  int_SFF_XXXX SFF_167 (bistsel,TDO_ISR,tdo_166,int_hold,g6601,CK,clockdr,updatedr,shiftdr,tdo_167,g25);
  int_SFF_XXXX SFF_168 (bistsel,TDO_ISR,tdo_167,int_hold,g5875,CK,clockdr,updatedr,shiftdr,tdo_168,g204);
  int_SFF_XXXX SFF_169 (bistsel,TDO_ISR,tdo_168,int_hold,g4425,CK,clockdr,updatedr,shiftdr,tdo_169,g658);
  int_SFF_XXXX SFF_170 (bistsel,TDO_ISR,tdo_169,int_hold,g5329,CK,clockdr,updatedr,shiftdr,tdo_170,g650);
  int_SFF_XXXX SFF_171 (bistsel,TDO_ISR,tdo_170,int_hold,g5695,CK,clockdr,updatedr,shiftdr,tdo_171,g378);
  int_SFF_XXXX SFF_172 (bistsel,TDO_ISR,tdo_171,int_hold,g6499,CK,clockdr,updatedr,shiftdr,tdo_172,g508);
  int_SFF_XXXX SFF_173 (bistsel,TDO_ISR,tdo_172,int_hold,g6825,CK,clockdr,updatedr,shiftdr,tdo_173,g548);
  int_SFF_XXXX SFF_174 (bistsel,TDO_ISR,tdo_173,int_hold,g5693,CK,clockdr,updatedr,shiftdr,tdo_174,g370);
  int_SFF_XXXX SFF_175 (bistsel,TDO_ISR,tdo_174,int_hold,g4850,CK,clockdr,updatedr,shiftdr,tdo_175,g406);
  int_SFF_XXXX SFF_176 (bistsel,TDO_ISR,tdo_175,int_hold,g3237,CK,clockdr,updatedr,shiftdr,tdo_176,g236);
  int_SFF_XXXX SFF_177 (bistsel,TDO_ISR,tdo_176,int_hold,g6497,CK,clockdr,updatedr,shiftdr,tdo_177,g500);
  int_SFF_XXXX SFF_178 (bistsel,TDO_ISR,tdo_177,int_hold,g6100,CK,clockdr,updatedr,shiftdr,tdo_178,g205);
  int_SFF_XXXX SFF_179 (bistsel,TDO_ISR,tdo_178,int_hold,g6509,CK,clockdr,updatedr,shiftdr,tdo_179,g197);
  int_SFF_XXXX SFF_180 (bistsel,TDO_ISR,tdo_179,int_hold,g4128,CK,clockdr,updatedr,shiftdr,tdo_180,g666);
  int_SFF_XXXX SFF_181 (bistsel,TDO_ISR,tdo_180,int_hold,g4116,CK,clockdr,updatedr,shiftdr,tdo_181,g114);
  int_SFF_XXXX SFF_182 (bistsel,TDO_ISR,tdo_181,int_hold,g6503,CK,clockdr,updatedr,shiftdr,tdo_182,g524);
  int_SFF_XXXX SFF_183 (bistsel,TDO_ISR,tdo_182,int_hold,g3241,CK,clockdr,updatedr,shiftdr,tdo_183,g260);
  int_SFF_XXXX SFF_184 (bistsel,TDO_ISR,tdo_183,int_hold,g6277,CK,clockdr,updatedr,shiftdr,tdo_184,g111);
  int_SFF_XXXX SFF_185 (bistsel,TDO_ISR,tdo_184,int_hold,g5139,CK,clockdr,updatedr,shiftdr,tdo_185,g131);
  int_SFF_XXXX SFF_186 (bistsel,TDO_ISR,tdo_185,int_hold,g6598,CK,clockdr,updatedr,shiftdr,tdo_186,g7);
  int_SFF_XXXX SFF_187 (bistsel,TDO_ISR,tdo_186,int_hold,g6600,CK,clockdr,updatedr,shiftdr,tdo_187,g19);
  int_SFF_XXXX SFF_188 (bistsel,TDO_ISR,tdo_187,int_hold,g4129,CK,clockdr,updatedr,shiftdr,tdo_188,g677);
  int_SFF_XXXX SFF_189 (bistsel,TDO_ISR,tdo_188,int_hold,g6593,CK,clockdr,updatedr,shiftdr,tdo_189,g582);
  int_SFF_XXXX SFF_190 (bistsel,TDO_ISR,tdo_189,int_hold,g6801,CK,clockdr,updatedr,shiftdr,tdo_190,g485);
  int_SFF_XXXX SFF_191 (bistsel,TDO_ISR,tdo_190,int_hold,g4426,CK,clockdr,updatedr,shiftdr,tdo_191,g699);
  int_SFF_XXXX SFF_192 (bistsel,TDO_ISR,tdo_191,int_hold,g5474,CK,clockdr,updatedr,shiftdr,tdo_192,g193);
  int_SFF_XXXX SFF_193 (bistsel,TDO_ISR,tdo_192,int_hold,g5140,CK,clockdr,updatedr,shiftdr,tdo_193,g135);
  int_SFF_XXXX SFF_194 (bistsel,TDO_ISR,tdo_193,int_hold,g5696,CK,clockdr,updatedr,shiftdr,tdo_194,g382);
  int_SFF_XXXX SFF_195 (bistsel,TDO_ISR,tdo_194,int_hold,g4852,CK,clockdr,updatedr,shiftdr,tdo_195,g414);
  int_SFF_XXXX SFF_196 (bistsel,TDO_ISR,tdo_195,int_hold,g4848,CK,clockdr,updatedr,shiftdr,tdo_196,g434);
  int_SFF_XXXX SFF_197 (bistsel,TDO_ISR,tdo_196,int_hold,g4659,CK,clockdr,updatedr,shiftdr,tdo_197,g266);
  int_SFF_XXXX SFF_198 (bistsel,TDO_ISR,tdo_197,int_hold,g6583,CK,clockdr,updatedr,shiftdr,tdo_198,g49);
  int_SFF_XXXX SFF_199 (bistsel,TDO_ISR,tdo_198,int_hold,g6402,CK,clockdr,updatedr,shiftdr,tdo_199,g152);
  int_SFF_XXXX SFF_200 (bistsel,TDO_ISR,tdo_199,int_hold,g4144,CK,clockdr,updatedr,shiftdr,tdo_200,g692);
  int_SFF_XXXX SFF_201 (bistsel,TDO_ISR,tdo_200,int_hold,g6104,CK,clockdr,updatedr,shiftdr,tdo_201,g277);
  int_SFF_XXXX SFF_202 (bistsel,TDO_ISR,tdo_201,int_hold,g6941,CK,clockdr,updatedr,shiftdr,tdo_202,g127);
  int_SFF_XXXX SFF_203 (bistsel,TDO_ISR,tdo_202,int_hold,g6403,CK,clockdr,updatedr,shiftdr,tdo_203,g161);
  int_SFF_XXXX SFF_204 (bistsel,TDO_ISR,tdo_203,int_hold,g6500,CK,clockdr,updatedr,shiftdr,tdo_204,g512);
  int_SFF_XXXX SFF_205 (bistsel,TDO_ISR,tdo_204,int_hold,g6508,CK,clockdr,updatedr,shiftdr,tdo_205,g532);
  int_SFF_XXXX SFF_206 (bistsel,TDO_ISR,tdo_205,int_hold,g6586,CK,clockdr,updatedr,shiftdr,tdo_206,g64);
  int_SFF_XXXX SFF_207 (bistsel,TDO_ISR,tdo_206,int_hold,g4146,CK,clockdr,updatedr,shiftdr,tdo_207,g694);
  int_SFF_XXXX SFF_208 (bistsel,TDO_ISR,tdo_207,int_hold,g4143,CK,clockdr,updatedr,shiftdr,tdo_208,g691);
  int_SFF_XXXX SFF_209 (bistsel,TDO_ISR,tdo_208,int_hold,g6720,CK,clockdr,updatedr,shiftdr,tdo_209,g1);
  int_SFF_XXXX SFF_210 (bistsel,TDO_ISR,tdo_209,int_hold,g6585,CK,clockdr,updatedr,shiftdr,TDO_ISR,g59);

  not NOT_0(I8854,g6696);
  not NOT_1(g1289,I2272);
  not NOT_2(I9125,g6855);
  not NOT_3(I6783,g4822);
  not NOT_4(I4424,g2097);
  not NOT_5(g6895,I9152);
  not NOT_6(g1835,I2919);
  not NOT_7(I3040,g1770);
  not NOT_8(g6837,g6822);
  not NOT_9(I7466,g5624);
  not NOT_10(I4809,g2974);
  not NOT_11(g3537,I4757);
  not NOT_12(g5457,g5304);
  not NOT_13(g6062,g5824);
  not NOT_14(g4040,I5343);
  not NOT_15(I6001,g4162);
  not NOT_16(g5549,g5331);
  not NOT_17(I4477,g3063);
  not NOT_18(g3612,I4809);
  not NOT_19(I7055,g5318);
  not NOT_20(g2892,g1982);
  not NOT_21(I5264,g3638);
  not NOT_22(I2225,g696);
  not NOT_23(g4123,I5451);
  not NOT_24(g4323,g4086);
  not NOT_25(g908,I1932);
  not NOT_26(I5933,g4346);
  not NOT_27(I8252,g6294);
  not NOT_28(I2473,g971);
  not NOT_29(I7333,g5386);
  not NOT_30(I8812,g6688);
  not NOT_31(g1674,g985);
  not NOT_32(I3528,g1422);
  not NOT_33(I8958,g6774);
  not NOT_34(I5050,g3246);
  not NOT_35(g3234,I4501);
  not NOT_36(I2324,g1209);
  not NOT_37(g2945,I4133);
  not NOT_38(g5121,I6775);
  not NOT_39(g1997,g1398);
  not NOT_40(g3128,I4375);
  not NOT_41(I8005,g6110);
  not NOT_42(g1541,g1094);
  not NOT_43(g5670,g5527);
  not NOT_44(g2738,g2327);
  not NOT_45(g6842,I9047);
  not NOT_46(g4528,I6096);
  not NOT_47(g2244,I3379);
  not NOT_48(g6192,g5946);
  not NOT_49(g2709,I3864);
  not NOT_50(g1332,I2349);
  not NOT_51(g4530,I6102);
  not NOT_52(g1680,g1011);
  not NOT_53(g2078,g1345);
  not NOT_54(g1209,I2215);
  not NOT_55(I3010,g1504);
  not NOT_56(g5813,I7612);
  not NOT_57(I7509,g5587);
  not NOT_58(I5379,g3940);
  not NOT_59(g3800,g3388);
  not NOT_60(g2907,g1914);
  not NOT_61(g6854,I9085);
  not NOT_62(g2035,I3144);
  not NOT_63(g2959,g1861);
  not NOT_64(g6941,I9236);
  not NOT_65(g4010,g3601);
  not NOT_66(I2287,g927);
  not NOT_67(I4273,g2197);
  not NOT_68(I8270,g6300);
  not NOT_69(g5740,I7501);
  not NOT_70(I5777,g3807);
  not NOT_71(g2876,g1943);
  not NOT_72(g873,g306);
  not NOT_73(g4839,I6525);
  not NOT_74(I5882,g3871);
  not NOT_75(g2656,I3800);
  not NOT_76(I8473,g6485);
  not NOT_77(I2199,g33);
  not NOT_78(g900,I1927);
  not NOT_79(g6708,I8834);
  not NOT_80(I2399,g729);
  not NOT_81(I3278,g1695);
  not NOT_82(g6520,I8476);
  not NOT_83(g940,g64);
  not NOT_84(I6677,g4757);
  not NOT_85(g3902,g3575);
  not NOT_86(g5687,g5567);
  not NOT_87(g2915,g1931);
  not NOT_88(g847,g590);
  not NOT_89(I3235,g1807);
  not NOT_90(I3343,g1623);
  not NOT_91(g6431,I8295);
  not NOT_92(g709,g114);
  not NOT_93(g6812,I8984);
  not NOT_94(I6576,g4700);
  not NOT_95(g749,I1847);
  not NOT_96(g3090,I4331);
  not NOT_97(I9107,g6855);
  not NOT_98(g2214,I3349);
  not NOT_99(g4618,g4246);
  not NOT_100(g6376,g6267);
  not NOT_101(g4143,I5511);
  not NOT_102(I6349,g4569);
  not NOT_103(g4343,g4011);
  not NOT_104(I5674,g4003);
  not NOT_105(I8177,g6173);
  not NOT_106(g2110,g1381);
  not NOT_107(I3134,g1336);
  not NOT_108(g6405,I8229);
  not NOT_109(I3334,g1330);
  not NOT_110(I7197,g5431);
  not NOT_111(g4566,g4198);
  not NOT_112(I7397,g5561);
  not NOT_113(I4534,g2858);
  not NOT_114(g1714,g1110);
  not NOT_115(I4961,g3597);
  not NOT_116(g2663,g2308);
  not NOT_117(g3456,g2640);
  not NOT_118(g5141,I6801);
  not NOT_119(g922,I1947);
  not NOT_120(g4693,I6283);
  not NOT_121(g4134,I5484);
  not NOT_122(g5570,g5392);
  not NOT_123(g5860,g5634);
  not NOT_124(g4334,g3733);
  not NOT_125(I3804,g2575);
  not NOT_126(I2207,g7);
  not NOT_127(I5153,g3330);
  not NOT_128(g3355,g3100);
  not NOT_129(g5645,g5537);
  not NOT_130(g6733,I8891);
  not NOT_131(g5691,g5568);
  not NOT_132(g4804,g4473);
  not NOT_133(I9047,g6838);
  not NOT_134(I4414,g2090);
  not NOT_135(g6610,I8696);
  not NOT_136(g2877,g2434);
  not NOT_137(I4903,g3223);
  not NOT_138(g6796,I8958);
  not NOT_139(g3063,I4288);
  not NOT_140(I3313,g1337);
  not NOT_141(g5879,g5770);
  not NOT_142(g3463,g2682);
  not NOT_143(I4513,g2765);
  not NOT_144(g1623,I2578);
  not NOT_145(g5358,I7012);
  not NOT_146(I3202,g1812);
  not NOT_147(I2215,g695);
  not NOT_148(g4113,I5421);
  not NOT_149(g1076,I2115);
  not NOT_150(g6069,g5791);
  not NOT_151(I7817,g5924);
  not NOT_152(g6540,g6474);
  not NOT_153(I6352,g4564);
  not NOT_154(I1865,g279);
  not NOT_155(g4202,I5622);
  not NOT_156(I6867,g5082);
  not NOT_157(I5511,g3876);
  not NOT_158(g5587,I7349);
  not NOT_159(I8144,g6182);
  not NOT_160(g1175,g42);
  not NOT_161(g1375,I2411);
  not NOT_162(g3118,I4366);
  not NOT_163(g3318,I4593);
  not NOT_164(g2464,I3596);
  not NOT_165(g3872,g3312);
  not NOT_166(g4494,I6004);
  not NOT_167(I2870,g1161);
  not NOT_168(g4518,I6066);
  not NOT_169(I4288,g2215);
  not NOT_170(g5615,I7372);
  not NOT_171(g4567,I6139);
  not NOT_172(I4382,g2265);
  not NOT_173(I3776,g2044);
  not NOT_174(g3057,I4282);
  not NOT_175(I5600,g3821);
  not NOT_176(I3593,g1295);
  not NOT_177(I2825,g1143);
  not NOT_178(g1285,g852);
  not NOT_179(g3457,g2653);
  not NOT_180(g5174,g5099);
  not NOT_181(I6386,g4462);
  not NOT_182(I3965,g2268);
  not NOT_183(I8488,g6426);
  not NOT_184(g6849,I9074);
  not NOT_185(I6599,g4823);
  not NOT_186(I2408,g719);
  not NOT_187(g3834,I5027);
  not NOT_188(g2295,g1578);
  not NOT_189(g1384,I2420);
  not NOT_190(g1339,I2370);
  not NOT_191(g5545,g5331);
  not NOT_192(I6170,g4343);
  not NOT_193(I9128,g6864);
  not NOT_194(g6898,I9161);
  not NOT_195(g1838,g1595);
  not NOT_196(g6900,I9167);
  not NOT_197(g2194,I3331);
  not NOT_198(g6797,I8961);
  not NOT_199(g2394,I3537);
  not NOT_200(I3050,g1439);
  not NOT_201(I3641,g1491);
  not NOT_202(I2943,g1715);
  not NOT_203(I5736,g4022);
  not NOT_204(g6510,I8450);
  not NOT_205(I6280,g4430);
  not NOT_206(g4933,I6625);
  not NOT_207(g5420,I7086);
  not NOT_208(g4521,I6075);
  not NOT_209(g1672,g1094);
  not NOT_210(I7058,g5281);
  not NOT_211(I2887,g1123);
  not NOT_212(I2122,g689);
  not NOT_213(g1477,g952);
  not NOT_214(g3232,I4495);
  not NOT_215(I2228,g15);
  not NOT_216(g5794,I7593);
  not NOT_217(g1643,I2608);
  not NOT_218(I4495,g3022);
  not NOT_219(I4437,g2108);
  not NOT_220(g2705,I3858);
  not NOT_221(g3813,g3258);
  not NOT_222(I8650,g6529);
  not NOT_223(I3379,g1647);
  not NOT_224(g2242,I3373);
  not NOT_225(g1205,g45);
  not NOT_226(I2033,g678);
  not NOT_227(I5871,g3744);
  not NOT_228(g774,I1859);
  not NOT_229(g6819,I8994);
  not NOT_230(g6694,I8800);
  not NOT_231(g4379,I5848);
  not NOT_232(g5905,g5852);
  not NOT_233(g3519,g2740);
  not NOT_234(I7856,g5994);
  not NOT_235(g921,g111);
  not NOT_236(g1551,g1011);
  not NOT_237(g1742,I2756);
  not NOT_238(I4752,g2859);
  not NOT_239(g6488,g6367);
  not NOT_240(g2254,I3391);
  not NOT_241(I8594,g6446);
  not NOT_242(g2814,I4023);
  not NOT_243(g4289,I5746);
  not NOT_244(g4658,I6247);
  not NOT_245(I6756,g4775);
  not NOT_246(g6701,I8821);
  not NOT_247(I8972,g6795);
  not NOT_248(I3271,g1748);
  not NOT_249(I2845,g1193);
  not NOT_250(g5300,I6952);
  not NOT_251(g2350,I3502);
  not NOT_252(I8806,g6686);
  not NOT_253(I3611,g1771);
  not NOT_254(I2137,g1);
  not NOT_255(I8943,g6774);
  not NOT_256(I2337,g1209);
  not NOT_257(I2913,g1792);
  not NOT_258(g1754,I2773);
  not NOT_259(g6886,I9125);
  not NOT_260(g2409,g1815);
  not NOT_261(g894,I1917);
  not NOT_262(g1273,g839);
  not NOT_263(I5424,g3725);
  not NOT_264(I6403,g4492);
  not NOT_265(g6314,I8044);
  not NOT_266(g4799,g4485);
  not NOT_267(I9155,g6882);
  not NOT_268(g2836,g2509);
  not NOT_269(g2212,I3343);
  not NOT_270(I6763,g4780);
  not NOT_271(g3860,I5081);
  not NOT_272(g2967,I4166);
  not NOT_273(g6825,I9008);
  not NOT_274(g5440,g5266);
  not NOT_275(g3710,g3029);
  not NOT_276(I5523,g3840);
  not NOT_277(g843,g574);
  not NOT_278(g1543,g1006);
  not NOT_279(g4132,I5478);
  not NOT_280(g6408,g6283);
  not NOT_281(g4153,I5545);
  not NOT_282(I6359,g4566);
  not NOT_283(g6136,I7856);
  not NOT_284(g2822,I4031);
  not NOT_285(I8891,g6706);
  not NOT_286(I8913,g6743);
  not NOT_287(I2692,g1037);
  not NOT_288(g6594,I8650);
  not NOT_289(g946,g361);
  not NOT_290(g1729,I2731);
  not NOT_291(I5551,g4059);
  not NOT_292(g4802,I6470);
  not NOT_293(g3962,I5214);
  not NOT_294(I2154,g14);
  not NOT_295(I4189,g2159);
  not NOT_296(I5499,g3847);
  not NOT_297(g5151,I6819);
  not NOT_298(g3158,I4398);
  not NOT_299(g6806,I8978);
  not NOT_300(I4706,g2877);
  not NOT_301(g5875,I7637);
  not NOT_302(g5530,I7270);
  not NOT_303(I9167,g6878);
  not NOT_304(I5926,g4153);
  not NOT_305(g2921,g1950);
  not NOT_306(g6065,g5784);
  not NOT_307(I6315,g4446);
  not NOT_308(I4371,g2555);
  not NOT_309(g6887,I9128);
  not NOT_310(I4429,g2102);
  not NOT_311(g6122,I7838);
  not NOT_312(g6465,I8329);
  not NOT_313(g6322,I8056);
  not NOT_314(g1660,g985);
  not NOT_315(g1946,I3053);
  not NOT_316(g6230,g6040);
  not NOT_317(g5010,I6646);
  not NOT_318(g4511,I6045);
  not NOT_319(I6874,g4861);
  not NOT_320(g2895,g1894);
  not NOT_321(g6033,g5824);
  not NOT_322(g2837,g2512);
  not NOT_323(I2979,g1263);
  not NOT_324(I3864,g2044);
  not NOT_325(g5884,g5864);
  not NOT_326(I8342,g6314);
  not NOT_327(I2218,g11);
  not NOT_328(g1513,g878);
  not NOT_329(I2312,g897);
  not NOT_330(I3714,g1852);
  not NOT_331(I4297,g2555);
  not NOT_332(I8255,g6292);
  not NOT_333(I8815,g6689);
  not NOT_334(g4492,I5998);
  not NOT_335(I1868,g280);
  not NOT_336(I7608,g5605);
  not NOT_337(I5862,g3863);
  not NOT_338(g1679,g985);
  not NOT_339(g1378,I2414);
  not NOT_340(g4714,I6324);
  not NOT_341(I2293,g971);
  not NOT_342(g5278,I6937);
  not NOT_343(g3284,g3019);
  not NOT_344(I4684,g2687);
  not NOT_345(I8497,g6481);
  not NOT_346(g3239,I4516);
  not NOT_347(I6537,g4711);
  not NOT_348(g3545,g3085);
  not NOT_349(g2788,I3983);
  not NOT_350(g6137,I7859);
  not NOT_351(g5667,g5524);
  not NOT_352(g6891,I9140);
  not NOT_353(g1831,I2907);
  not NOT_354(g1335,I2358);
  not NOT_355(g3380,g2831);
  not NOT_356(I4791,g2814);
  not NOT_357(g6337,I8089);
  not NOT_358(I4309,g2525);
  not NOT_359(I2828,g1193);
  not NOT_360(g3832,I5023);
  not NOT_361(g1288,I2269);
  not NOT_362(g5566,I7318);
  not NOT_363(g3853,I5068);
  not NOT_364(I3736,g2460);
  not NOT_365(I6612,g4660);
  not NOT_366(I7161,g5465);
  not NOT_367(I7361,g5566);
  not NOT_368(g2842,I4050);
  not NOT_369(g1805,I2854);
  not NOT_370(I6417,g4617);
  not NOT_371(I3623,g1491);
  not NOT_372(g4262,I5713);
  not NOT_373(I7051,g5219);
  not NOT_374(I2221,g43);
  not NOT_375(g3559,g2603);
  not NOT_376(g4736,I6366);
  not NOT_377(g2485,I3614);
  not NOT_378(I7451,g5597);
  not NOT_379(I2703,g1189);
  not NOT_380(I8267,g6297);
  not NOT_381(g4623,g4262);
  not NOT_382(g1947,I3056);
  not NOT_383(I5885,g3746);
  not NOT_384(I7999,g6137);
  not NOT_385(g878,g639);
  not NOT_386(I7146,g5231);
  not NOT_387(I6330,g4560);
  not NOT_388(I7346,g5531);
  not NOT_389(I3871,g2145);
  not NOT_390(I8329,g6305);
  not NOT_391(g4375,I5840);
  not NOT_392(g4871,I6599);
  not NOT_393(I8761,g6563);
  not NOT_394(g3204,I4441);
  not NOT_395(g4722,I6346);
  not NOT_396(g710,g128);
  not NOT_397(I4498,g2686);
  not NOT_398(g829,g323);
  not NOT_399(g5113,I6753);
  not NOT_400(g1632,g760);
  not NOT_401(g1037,I2067);
  not NOT_402(g3100,I4347);
  not NOT_403(I8828,g6661);
  not NOT_404(g6726,I8872);
  not NOT_405(g6497,I8411);
  not NOT_406(g1653,I2630);
  not NOT_407(g2640,I3782);
  not NOT_408(I8727,g6536);
  not NOT_409(g2031,I3140);
  not NOT_410(I5436,g3729);
  not NOT_411(g2252,I3385);
  not NOT_412(g5908,g5753);
  not NOT_413(g2958,g1861);
  not NOT_414(I7472,g5626);
  not NOT_415(g2176,I3319);
  not NOT_416(I2716,g1115);
  not NOT_417(I5831,g3842);
  not NOT_418(I2349,g1160);
  not NOT_419(g4139,I5499);
  not NOT_420(I5182,g3271);
  not NOT_421(g5518,I7258);
  not NOT_422(g5567,g5418);
  not NOT_423(I5382,g3952);
  not NOT_424(g2405,I3543);
  not NOT_425(I2848,g1193);
  not NOT_426(g1917,I3016);
  not NOT_427(g2829,g2491);
  not NOT_428(g2765,I3946);
  not NOT_429(I7116,g5299);
  not NOT_430(I4019,g1841);
  not NOT_431(g4424,I5923);
  not NOT_432(I6090,g4393);
  not NOT_433(I4362,g2555);
  not NOT_434(I3672,g1656);
  not NOT_435(g3040,I4255);
  not NOT_436(I3077,g1439);
  not NOT_437(g4809,I6485);
  not NOT_438(g5593,I7355);
  not NOT_439(g3440,I4678);
  not NOT_440(g3969,I5233);
  not NOT_441(g6312,I8040);
  not NOT_442(I6366,g4569);
  not NOT_443(I4452,g2117);
  not NOT_444(g2974,I4173);
  not NOT_445(g6401,I8217);
  not NOT_446(g895,g139);
  not NOT_447(I6456,g4633);
  not NOT_448(g4523,I6081);
  not NOT_449(g1233,I2231);
  not NOT_450(I6649,g4693);
  not NOT_451(g4643,g4293);
  not NOT_452(g5264,g4943);
  not NOT_453(I9158,g6887);
  not NOT_454(g1054,g485);
  not NOT_455(g5160,g5099);
  not NOT_456(g2796,I3999);
  not NOT_457(I6355,g4569);
  not NOT_458(g2473,I3605);
  not NOT_459(I3099,g1519);
  not NOT_460(I8576,g6436);
  not NOT_461(g1770,I2805);
  not NOT_462(I8866,g6701);
  not NOT_463(I3304,g1740);
  not NOT_464(I4486,g3093);
  not NOT_465(g5521,I7261);
  not NOT_466(I3499,g1450);
  not NOT_467(I8716,g6518);
  not NOT_468(g1725,g1113);
  not NOT_469(I7596,g5605);
  not NOT_470(g6727,I8875);
  not NOT_471(g3875,I5106);
  not NOT_472(g2324,I3478);
  not NOT_473(I4504,g2726);
  not NOT_474(I2119,g688);
  not NOT_475(g5450,g5292);
  not NOT_476(I5037,g3705);
  not NOT_477(g5996,g5824);
  not NOT_478(g4104,I5394);
  not NOT_479(g6592,I8644);
  not NOT_480(g4099,I5379);
  not NOT_481(g4499,I6015);
  not NOT_482(I2352,g1161);
  not NOT_483(I6063,g4381);
  not NOT_484(g6746,I8916);
  not NOT_485(I2867,g1143);
  not NOT_486(I8699,g6573);
  not NOT_487(g2177,I3322);
  not NOT_488(g5179,g5099);
  not NOT_489(g5379,I7035);
  not NOT_490(I2893,g1236);
  not NOT_491(g5878,I7646);
  not NOT_492(I3044,g1257);
  not NOT_493(g1189,I2196);
  not NOT_494(g3839,I5040);
  not NOT_495(g6932,I9217);
  not NOT_496(g4273,I5728);
  not NOT_497(g5658,g5512);
  not NOT_498(g6624,I8730);
  not NOT_499(I6118,g4406);
  not NOT_500(I6318,g4447);
  not NOT_501(I3983,g2276);
  not NOT_502(g2849,g2577);
  not NOT_503(I3572,g1295);
  not NOT_504(g1787,I2835);
  not NOT_505(I5442,g3731);
  not NOT_506(I4678,g2670);
  not NOT_507(I6057,g4379);
  not NOT_508(I8524,g6496);
  not NOT_509(I4331,g2555);
  not NOT_510(I8644,g6526);
  not NOT_511(I3543,g1461);
  not NOT_512(I6989,g5307);
  not NOT_513(I2614,g1123);
  not NOT_514(g1675,g1101);
  not NOT_515(I2370,g1123);
  not NOT_516(I2125,g698);
  not NOT_517(g3235,I4504);
  not NOT_518(g3343,g3090);
  not NOT_519(I5233,g3571);
  not NOT_520(I2821,g1221);
  not NOT_521(g4712,I6318);
  not NOT_522(g985,g638);
  not NOT_523(g6576,g6487);
  not NOT_524(I6549,g4699);
  not NOT_525(I8258,g6293);
  not NOT_526(I8818,g6690);
  not NOT_527(I3534,g1295);
  not NOT_528(g2245,I3382);
  not NOT_529(I3729,g2436);
  not NOT_530(I3961,g1835);
  not NOT_531(I5454,g3874);
  not NOT_532(g2291,I3434);
  not NOT_533(g5997,g5854);
  not NOT_534(g4534,I6114);
  not NOT_535(I3927,g2245);
  not NOT_536(I5532,g3861);
  not NOT_537(g1684,I2668);
  not NOT_538(g6699,I8815);
  not NOT_539(g1639,g815);
  not NOT_540(g1338,I2367);
  not NOT_541(g1963,I3074);
  not NOT_542(I8186,g6179);
  not NOT_543(I6321,g4559);
  not NOT_544(I4226,g2525);
  not NOT_545(g1109,I2137);
  not NOT_546(g1791,I2845);
  not NOT_547(I8975,g6791);
  not NOT_548(I3946,g2256);
  not NOT_549(g889,g310);
  not NOT_550(I2306,g896);
  not NOT_551(g3792,g3388);
  not NOT_552(I6625,g4745);
  not NOT_553(g2819,g2467);
  not NOT_554(g4014,I5316);
  not NOT_555(I8426,g6424);
  not NOT_556(I5412,g4034);
  not NOT_557(g4660,I6253);
  not NOT_558(I6253,g4608);
  not NOT_559(g2088,I3202);
  not NOT_560(g2923,g1969);
  not NOT_561(I4173,g2408);
  not NOT_562(I8614,g6537);
  not NOT_563(I3513,g1450);
  not NOT_564(g2488,I3617);
  not NOT_565(g1759,I2782);
  not NOT_566(I2756,g1175);
  not NOT_567(g2701,I3855);
  not NOT_568(I7190,g5432);
  not NOT_569(I8821,g6691);
  not NOT_570(g6524,I8488);
  not NOT_571(I6740,g4781);
  not NOT_572(g4513,I6051);
  not NOT_573(I8984,g6794);
  not NOT_574(I7501,g5596);
  not NOT_575(g1957,I3068);
  not NOT_576(g2215,I3352);
  not NOT_577(g6119,I7829);
  not NOT_578(I2904,g1256);
  not NOT_579(g6319,I8051);
  not NOT_580(g1049,g266);
  not NOT_581(g5901,g5753);
  not NOT_582(g2886,g1966);
  not NOT_583(I6552,g4702);
  not NOT_584(I4059,g1878);
  not NOT_585(g4036,I5337);
  not NOT_586(g3094,I4337);
  not NOT_587(I4459,g2134);
  not NOT_588(I8544,g6453);
  not NOT_589(g4679,I6269);
  not NOT_590(g6352,I8110);
  not NOT_591(g6818,I8991);
  not NOT_592(g6577,g6488);
  not NOT_593(I1847,g209);
  not NOT_594(I3288,g1710);
  not NOT_595(g3567,g3074);
  not NOT_596(I3382,g1284);
  not NOT_597(g1715,I2716);
  not NOT_598(g4135,I5487);
  not NOT_599(I7704,g5723);
  not NOT_600(g848,g594);
  not NOT_601(g5092,g4753);
  not NOT_602(g1498,I2479);
  not NOT_603(I2763,g1236);
  not NOT_604(g2870,g2296);
  not NOT_605(I3022,g1426);
  not NOT_606(I4261,g1857);
  not NOT_607(I2391,g774);
  not NOT_608(g4382,I5857);
  not NOT_609(g3776,g3466);
  not NOT_610(g6893,I9146);
  not NOT_611(g1833,I2913);
  not NOT_612(I3422,g1641);
  not NOT_613(g5574,g5407);
  not NOT_614(I3749,g2484);
  not NOT_615(g3593,g2997);
  not NOT_616(g6211,g5992);
  not NOT_617(g2650,I3794);
  not NOT_618(g5714,I7475);
  not NOT_619(g932,g337);
  not NOT_620(I8061,g6113);
  not NOT_621(g4805,g4473);
  not NOT_622(g4022,I5328);
  not NOT_623(g1584,g743);
  not NOT_624(g4422,g4111);
  not NOT_625(g6599,I8665);
  not NOT_626(g1539,g878);
  not NOT_627(I5109,g3710);
  not NOT_628(g2408,I3546);
  not NOT_629(I2159,g465);
  not NOT_630(I6570,g4719);
  not NOT_631(g2136,g1395);
  not NOT_632(I4664,g2924);
  not NOT_633(I8027,g6237);
  not NOT_634(I4246,g2194);
  not NOT_635(g2336,I3488);
  not NOT_636(g5580,I7336);
  not NOT_637(g716,I1832);
  not NOT_638(I3560,g1673);
  not NOT_639(g736,I1841);
  not NOT_640(I6525,g4770);
  not NOT_641(g2768,g2367);
  not NOT_642(g6370,I8174);
  not NOT_643(g2594,I3723);
  not NOT_644(g4798,I6464);
  not NOT_645(g6325,I8061);
  not NOT_646(g6821,g6785);
  not NOT_647(g4560,g4188);
  not NOT_648(g2806,g2446);
  not NOT_649(I3632,g1295);
  not NOT_650(g3450,I4688);
  not NOT_651(I3037,g1769);
  not NOT_652(g6939,I9230);
  not NOT_653(g1052,g668);
  not NOT_654(I3653,g1305);
  not NOT_655(I3102,g1426);
  not NOT_656(I2115,g687);
  not NOT_657(I2315,g1222);
  not NOT_658(I2811,g1209);
  not NOT_659(g6083,g5809);
  not NOT_660(g2887,g1858);
  not NOT_661(I2047,g682);
  not NOT_662(g6544,I8544);
  not NOT_663(I6607,g4745);
  not NOT_664(g4632,g4281);
  not NOT_665(g5889,g5742);
  not NOT_666(g5476,I7164);
  not NOT_667(g2934,g2004);
  not NOT_668(g2230,I3355);
  not NOT_669(g4437,I5948);
  not NOT_670(g4102,I5388);
  not NOT_671(g4302,g4068);
  not NOT_672(I5865,g3743);
  not NOT_673(g6106,I7814);
  not NOT_674(g4579,g4206);
  not NOT_675(g4869,g4662);
  not NOT_676(g6306,I8030);
  not NOT_677(I3752,g2044);
  not NOT_678(g5375,I7029);
  not NOT_679(I8107,g6136);
  not NOT_680(g4719,I6337);
  not NOT_681(g1730,g1114);
  not NOT_682(g3289,g3034);
  not NOT_683(g1504,I2485);
  not NOT_684(g3777,g3388);
  not NOT_685(I6587,g4803);
  not NOT_686(I8159,g6167);
  not NOT_687(I6111,g4404);
  not NOT_688(g3835,I5030);
  not NOT_689(I6311,g4444);
  not NOT_690(I8223,g6325);
  not NOT_691(g2096,I3212);
  not NOT_692(I9143,g6886);
  not NOT_693(g3882,I5119);
  not NOT_694(g1070,g94);
  not NOT_695(g2550,I3665);
  not NOT_696(I6615,g4745);
  not NOT_697(g3271,g3042);
  not NOT_698(I4671,g2928);
  not NOT_699(I2880,g1143);
  not NOT_700(g2845,g2565);
  not NOT_701(g1897,I2992);
  not NOT_702(g6622,I8724);
  not NOT_703(I2537,g971);
  not NOT_704(I5896,g3879);
  not NOT_705(g2195,I3334);
  not NOT_706(g4265,I5716);
  not NOT_707(g2891,g1884);
  not NOT_708(g2913,g1925);
  not NOT_709(g5139,I6795);
  not NOT_710(I3364,g1648);
  not NOT_711(g5384,g5220);
  not NOT_712(I9134,g6864);
  not NOT_713(I2272,g908);
  not NOT_714(g6904,I9179);
  not NOT_715(g4786,I6448);
  not NOT_716(g3799,g3388);
  not NOT_717(g6514,I8462);
  not NOT_718(g4364,I5825);
  not NOT_719(I8447,g6410);
  not NOT_720(I3770,g2145);
  not NOT_721(I5019,g3318);
  not NOT_722(I2417,g774);
  not NOT_723(g6403,I8223);
  not NOT_724(g5809,I7608);
  not NOT_725(I7683,g5702);
  not NOT_726(g6841,I9044);
  not NOT_727(g3541,g2643);
  not NOT_728(I2982,g1426);
  not NOT_729(g1678,I2658);
  not NOT_730(g4770,I6414);
  not NOT_731(g1006,I2047);
  not NOT_732(I2234,g697);
  not NOT_733(g1331,I2346);
  not NOT_734(g4296,I5753);
  not NOT_735(I2128,g18);
  not NOT_736(g3238,I4513);
  not NOT_737(I3553,g1305);
  not NOT_738(I6020,g4176);
  not NOT_739(g3332,g3079);
  not NOT_740(g5477,I7167);
  not NOT_741(I6420,g4618);
  not NOT_742(g6695,I8803);
  not NOT_743(I2330,g1122);
  not NOT_744(g3209,I4452);
  not NOT_745(I6507,g4644);
  not NOT_746(g4532,I6108);
  not NOT_747(g1682,g829);
  not NOT_748(g6107,I7817);
  not NOT_749(I9113,g6855);
  not NOT_750(I1856,g204);
  not NOT_751(g1305,I2293);
  not NOT_752(g6536,I8524);
  not NOT_753(g3802,g3388);
  not NOT_754(I5728,g4022);
  not NOT_755(g2481,I3608);
  not NOT_756(I7475,g5627);
  not NOT_757(g931,g54);
  not NOT_758(g1748,I2763);
  not NOT_759(g2692,I3840);
  not NOT_760(I4217,g2163);
  not NOT_761(g2097,I3215);
  not NOT_762(I4066,g2582);
  not NOT_763(g5551,I7295);
  not NOT_764(g5742,g5686);
  not NOT_765(g2726,I3886);
  not NOT_766(g5099,I6737);
  not NOT_767(g2497,I3626);
  not NOT_768(I5385,g3962);
  not NOT_769(g5304,I6956);
  not NOT_770(g2154,I3271);
  not NOT_771(g1755,I2776);
  not NOT_772(g4189,I5597);
  not NOT_773(I8978,g6792);
  not NOT_774(g4706,I6308);
  not NOT_775(g6416,I8258);
  not NOT_776(I8243,g6286);
  not NOT_777(I8417,g6420);
  not NOT_778(g3901,g3575);
  not NOT_779(I6630,g4745);
  not NOT_780(I7646,g5774);
  not NOT_781(I3675,g1491);
  not NOT_782(g6522,I8482);
  not NOT_783(g6115,g5879);
  not NOT_784(g1045,g699);
  not NOT_785(I3281,g1761);
  not NOT_786(I7039,g5309);
  not NOT_787(I7484,g5630);
  not NOT_788(g1173,I2185);
  not NOT_789(I4455,g2118);
  not NOT_790(I8629,g6544);
  not NOT_791(g5273,I6930);
  not NOT_792(I4133,g2040);
  not NOT_793(g1491,I2476);
  not NOT_794(g760,I1853);
  not NOT_795(g2783,I3979);
  not NOT_796(g4281,I5736);
  not NOT_797(g3600,I4791);
  not NOT_798(g2112,I3240);
  not NOT_799(g1283,g853);
  not NOT_800(g2312,I3462);
  not NOT_801(g1369,I2405);
  not NOT_802(I6750,g4771);
  not NOT_803(g6654,I8758);
  not NOT_804(g3714,g3041);
  not NOT_805(I7583,g5605);
  not NOT_806(I3684,g1733);
  not NOT_807(I5006,g3604);
  not NOT_808(I8800,g6684);
  not NOT_809(g1059,g702);
  not NOT_810(g1578,I2552);
  not NOT_811(g2001,I3112);
  not NOT_812(I5406,g3976);
  not NOT_813(g5572,g5399);
  not NOT_814(I3109,g1504);
  not NOT_815(I3791,g2044);
  not NOT_816(g2293,g1567);
  not NOT_817(g6880,I9107);
  not NOT_818(g6595,I8653);
  not NOT_819(g4138,I5496);
  not NOT_820(g1535,g1088);
  not NOT_821(g4639,g4289);
  not NOT_822(g6537,I8527);
  not NOT_823(g5543,g5331);
  not NOT_824(I3808,g2125);
  not NOT_825(I7276,g5375);
  not NOT_826(I5487,g3881);
  not NOT_827(I2355,g1177);
  not NOT_828(g4109,I5409);
  not NOT_829(g4309,g4074);
  not NOT_830(g2828,g2488);
  not NOT_831(g2830,g2494);
  not NOT_832(g2727,g2324);
  not NOT_833(g4808,g4473);
  not NOT_834(I2964,g1257);
  not NOT_835(g821,I1880);
  not NOT_836(g6612,I8702);
  not NOT_837(g5534,I7276);
  not NOT_838(g5729,I7494);
  not NOT_839(I6666,g4740);
  not NOT_840(I9179,g6875);
  not NOT_841(g1415,g1246);
  not NOT_842(g4707,I6311);
  not NOT_843(g6417,I8261);
  not NOT_844(I7404,g5541);
  not NOT_845(g3076,I4309);
  not NOT_846(I8512,g6441);
  not NOT_847(g3889,g3575);
  not NOT_848(I6528,g4815);
  not NOT_849(g1664,I2643);
  not NOT_850(g1246,I2237);
  not NOT_851(g6234,g6057);
  not NOT_852(I3575,g1305);
  not NOT_853(g5885,g5865);
  not NOT_854(g6328,I8066);
  not NOT_855(g1203,I2207);
  not NOT_856(I5445,g4040);
  not NOT_857(g5946,g5729);
  not NOT_858(g6542,I8538);
  not NOT_859(g6330,I8070);
  not NOT_860(g1721,I2721);
  not NOT_861(I5091,g3242);
  not NOT_862(I8056,g6109);
  not NOT_863(g2932,g1998);
  not NOT_864(I8456,g6417);
  not NOT_865(g5903,g5753);
  not NOT_866(I3833,g2266);
  not NOT_867(I2318,g1236);
  not NOT_868(g4715,I6327);
  not NOT_869(I2367,g1161);
  not NOT_870(I1924,g663);
  not NOT_871(g6800,I8966);
  not NOT_872(I5169,g3593);
  not NOT_873(I6410,g4473);
  not NOT_874(g4098,I5376);
  not NOT_875(g3500,g2647);
  not NOT_876(g4498,I6012);
  not NOT_877(I2057,g685);
  not NOT_878(g1502,g709);
  not NOT_879(I5059,g3259);
  not NOT_880(I5920,g4228);
  not NOT_881(I2457,g1253);
  not NOT_882(I3584,g1678);
  not NOT_883(I5868,g3864);
  not NOT_884(I2989,g1519);
  not NOT_885(I2193,g693);
  not NOT_886(g5436,I7116);
  not NOT_887(g3384,g2834);
  not NOT_888(g1940,I3047);
  not NOT_889(g2576,I3687);
  not NOT_890(g2866,g1905);
  not NOT_891(g5135,I6783);
  not NOT_892(g2716,I3871);
  not NOT_893(g3838,I5037);
  not NOT_894(I7906,g5912);
  not NOT_895(I3268,g1656);
  not NOT_896(I3019,g1755);
  not NOT_897(g3424,I4671);
  not NOT_898(g5382,I7042);
  not NOT_899(I5793,g3803);
  not NOT_900(I3419,g1287);
  not NOT_901(g6902,I9173);
  not NOT_902(I6143,g4237);
  not NOT_903(I6343,g4458);
  not NOT_904(g846,g586);
  not NOT_905(g1671,g985);
  not NOT_906(g5805,I7604);
  not NOT_907(I5415,g3723);
  not NOT_908(g6512,I8456);
  not NOT_909(I3452,g1450);
  not NOT_910(g4162,I5562);
  not NOT_911(g5022,I6666);
  not NOT_912(g1030,I2057);
  not NOT_913(I8279,g6307);
  not NOT_914(g3231,I4492);
  not NOT_915(g6490,g6371);
  not NOT_916(I2321,g898);
  not NOT_917(g6823,I9002);
  not NOT_918(g3477,g2692);
  not NOT_919(g6166,I7892);
  not NOT_920(g6366,I8162);
  not NOT_921(I6334,g4454);
  not NOT_922(I8872,g6695);
  not NOT_923(g2241,I3370);
  not NOT_924(g1564,g1030);
  not NOT_925(I7892,g5916);
  not NOT_926(I3086,g1439);
  not NOT_927(g6529,I8503);
  not NOT_928(I8843,g6658);
  not NOT_929(g6649,I8745);
  not NOT_930(I6555,g4703);
  not NOT_931(g1741,I2753);
  not NOT_932(I6792,g5097);
  not NOT_933(g3104,I4351);
  not NOT_934(I3385,g1318);
  not NOT_935(g2524,I3647);
  not NOT_936(g2644,I3788);
  not NOT_937(I8834,g6661);
  not NOT_938(g6698,I8812);
  not NOT_939(g1638,g754);
  not NOT_940(g839,g567);
  not NOT_941(I6621,g4745);
  not NOT_942(g2119,g1391);
  not NOT_943(I5502,g3853);
  not NOT_944(g1108,I2134);
  not NOT_945(I3025,g1439);
  not NOT_946(I2552,g971);
  not NOT_947(g5437,I7119);
  not NOT_948(g4385,I5862);
  not NOT_949(I3425,g1274);
  not NOT_950(I9092,g6855);
  not NOT_951(I4441,g2109);
  not NOT_952(g2818,g2464);
  not NOT_953(g2867,g1908);
  not NOT_954(g1883,g1797);
  not NOT_955(g5579,I7333);
  not NOT_956(I7478,g5628);
  not NOT_957(g4425,I5926);
  not NOT_958(I7035,g5150);
  not NOT_959(I5388,g3969);
  not NOT_960(I7517,g5593);
  not NOT_961(g2893,g1985);
  not NOT_962(g5752,I7509);
  not NOT_963(I8232,g6332);
  not NOT_964(g5917,I7683);
  not NOT_965(I6567,g4715);
  not NOT_966(g6720,I8854);
  not NOT_967(I3678,g1690);
  not NOT_968(g2975,I4176);
  not NOT_969(I5030,g3242);
  not NOT_970(I3331,g1631);
  not NOT_971(g1861,I2967);
  not NOT_972(g6367,I8165);
  not NOT_973(g1048,g492);
  not NOT_974(I5430,g3727);
  not NOT_975(g2599,I3729);
  not NOT_976(g5042,I6672);
  not NOT_977(g1711,I2712);
  not NOT_978(I3635,g1305);
  not NOT_979(g6652,I8752);
  not NOT_980(g5442,g5270);
  not NOT_981(g1055,g269);
  not NOT_982(I2570,g1222);
  not NOT_983(I2860,g1177);
  not NOT_984(g6057,g5824);
  not NOT_985(g4131,I5475);
  not NOT_986(I4743,g2594);
  not NOT_987(I3105,g1439);
  not NOT_988(g2170,I3301);
  not NOT_989(g2370,I3522);
  not NOT_990(g4406,I5913);
  not NOT_991(g6193,g5957);
  not NOT_992(g1333,I2352);
  not NOT_993(g2125,I3255);
  not NOT_994(I8552,g6455);
  not NOT_995(g1774,I2817);
  not NOT_996(g4766,I6406);
  not NOT_997(g4105,I5397);
  not NOT_998(g1846,I2940);
  not NOT_999(g5054,g4816);
  not NOT_1000(g4801,g4487);
  not NOT_1001(g6834,g6821);
  not NOT_1002(g4487,I5991);
  not NOT_1003(I7110,g5291);
  not NOT_1004(g3534,I4752);
  not NOT_1005(I5910,g3750);
  not NOT_1006(g5770,g5645);
  not NOT_1007(I3755,g2125);
  not NOT_1008(g5296,I6946);
  not NOT_1009(I8687,g6568);
  not NOT_1010(I6933,g5124);
  not NOT_1011(g2544,I3662);
  not NOT_1012(g6598,I8662);
  not NOT_1013(I5609,g3893);
  not NOT_1014(I4474,g3052);
  not NOT_1015(I2358,g1176);
  not NOT_1016(g3014,I4217);
  not NOT_1017(g6121,I7835);
  not NOT_1018(I7002,g5308);
  not NOT_1019(g766,I1856);
  not NOT_1020(g3885,I5124);
  not NOT_1021(g4226,g4050);
  not NOT_1022(g2106,g1378);
  not NOT_1023(g2306,g1743);
  not NOT_1024(I3373,g1320);
  not NOT_1025(g2790,g2413);
  not NOT_1026(g6232,g6048);
  not NOT_1027(I5217,g3673);
  not NOT_1028(I8570,g6433);
  not NOT_1029(I8860,g6699);
  not NOT_1030(I4480,g3073);
  not NOT_1031(g1994,I3105);
  not NOT_1032(g1290,I2275);
  not NOT_1033(I2275,g909);
  not NOT_1034(g6938,I9227);
  not NOT_1035(I5466,g3787);
  not NOT_1036(g4173,I5577);
  not NOT_1037(I8710,g6517);
  not NOT_1038(g2461,I3593);
  not NOT_1039(I7590,g5605);
  not NOT_1040(I3602,g1491);
  not NOT_1041(I3007,g1439);
  not NOT_1042(g2756,g2353);
  not NOT_1043(g2622,I3764);
  not NOT_1044(I3059,g1519);
  not NOT_1045(I3578,g1484);
  not NOT_1046(I3868,g2125);
  not NOT_1047(g5888,g5731);
  not NOT_1048(g1256,g838);
  not NOT_1049(g6519,I8473);
  not NOT_1050(I6289,g4433);
  not NOT_1051(I9024,g6803);
  not NOT_1052(I5448,g3960);
  not NOT_1053(I3767,g2125);
  not NOT_1054(g5787,g5685);
  not NOT_1055(g2904,g1991);
  not NOT_1056(g6552,I8552);
  not NOT_1057(g6606,I8684);
  not NOT_1058(g2446,I3581);
  not NOT_1059(I5333,g3491);
  not NOT_1060(I2284,g922);
  not NOT_1061(g1381,I2417);
  not NOT_1062(g4718,I6334);
  not NOT_1063(g4767,g4601);
  not NOT_1064(I3261,g1783);
  not NOT_1065(g1847,I2943);
  not NOT_1066(I4688,g3207);
  not NOT_1067(I5774,g3807);
  not NOT_1068(I9077,g6845);
  not NOT_1069(I8659,g6523);
  not NOT_1070(g4535,g4173);
  not NOT_1071(I4976,g3575);
  not NOT_1072(g1685,I2671);
  not NOT_1073(g2145,I3268);
  not NOT_1074(I8506,g6483);
  not NOT_1075(g2841,g2541);
  not NOT_1076(g4582,g4210);
  not NOT_1077(g3022,I4229);
  not NOT_1078(g2391,I3534);
  not NOT_1079(g6586,I8626);
  not NOT_1080(g952,I2029);
  not NOT_1081(g1263,g846);
  not NOT_1082(g964,g357);
  not NOT_1083(I2420,g791);
  not NOT_1084(g2695,I3843);
  not NOT_1085(g2637,I3779);
  not NOT_1086(g1950,I3059);
  not NOT_1087(g5138,I6792);
  not NOT_1088(g4227,g4059);
  not NOT_1089(I7295,g5439);
  not NOT_1090(g5791,I7590);
  not NOT_1091(g3798,g3388);
  not NOT_1092(I9104,g6864);
  not NOT_1093(g5309,g5063);
  not NOT_1094(g2159,I3284);
  not NOT_1095(g6570,I8594);
  not NOT_1096(g4246,I5692);
  not NOT_1097(I6132,g4219);
  not NOT_1098(I8174,g6173);
  not NOT_1099(g6525,I8491);
  not NOT_1100(g6710,I8840);
  not NOT_1101(I5418,g4036);
  not NOT_1102(I6680,g4713);
  not NOT_1103(g4721,I6343);
  not NOT_1104(g1631,I2588);
  not NOT_1105(g2416,I3556);
  not NOT_1106(g3095,I4340);
  not NOT_1107(g3037,I4252);
  not NOT_1108(I3502,g1295);
  not NOT_1109(g1257,g845);
  not NOT_1110(g1101,I2125);
  not NOT_1111(I2204,g694);
  not NOT_1112(I2630,g1143);
  not NOT_1113(I5493,g3834);
  not NOT_1114(I8180,g6176);
  not NOT_1115(I4220,g2164);
  not NOT_1116(I7966,g6166);
  not NOT_1117(I8591,g6448);
  not NOT_1118(g2315,I3465);
  not NOT_1119(g5957,g5866);
  not NOT_1120(g6879,I9104);
  not NOT_1121(g6607,I8687);
  not NOT_1122(I6558,g4705);
  not NOT_1123(g4502,I6020);
  not NOT_1124(g5049,I6685);
  not NOT_1125(I9044,g6836);
  not NOT_1126(g927,I1958);
  not NOT_1127(I1942,g664);
  not NOT_1128(I4023,g2315);
  not NOT_1129(g3719,g3053);
  not NOT_1130(g6506,I8438);
  not NOT_1131(g5575,g5411);
  not NOT_1132(I8420,g6422);
  not NOT_1133(I3388,g1324);
  not NOT_1134(g2874,g1849);
  not NOT_1135(g3752,I4935);
  not NOT_1136(I5397,g3932);
  not NOT_1137(I3028,g1504);
  not NOT_1138(g4188,I5594);
  not NOT_1139(g6587,I8629);
  not NOT_1140(g4388,I5871);
  not NOT_1141(I5421,g3724);
  not NOT_1142(I3428,g1825);
  not NOT_1143(I2973,g1687);
  not NOT_1144(I7254,g5458);
  not NOT_1145(I7814,g5922);
  not NOT_1146(I3247,g1791);
  not NOT_1147(g3042,I4261);
  not NOT_1148(g6615,I8707);
  not NOT_1149(I7150,g5355);
  not NOT_1150(I4327,g2525);
  not NOT_1151(g4428,I5933);
  not NOT_1152(g3786,g3388);
  not NOT_1153(g5584,I7346);
  not NOT_1154(g5539,g5331);
  not NOT_1155(g5896,g5753);
  not NOT_1156(g1673,I2653);
  not NOT_1157(g6374,I8186);
  not NOT_1158(I3826,g2145);
  not NOT_1159(g3364,g3114);
  not NOT_1160(g3233,I4498);
  not NOT_1161(I8515,g6492);
  not NOT_1162(g4564,g4192);
  not NOT_1163(g3054,I4279);
  not NOT_1164(I5562,g4002);
  not NOT_1165(I4303,g1897);
  not NOT_1166(g2612,I3752);
  not NOT_1167(I8300,g6299);
  not NOT_1168(g6284,I8002);
  not NOT_1169(g2243,I3376);
  not NOT_1170(g3770,I4961);
  not NOT_1171(I9014,g6820);
  not NOT_1172(I3638,g1484);
  not NOT_1173(g1772,I2811);
  not NOT_1174(I5723,g3942);
  not NOT_1175(g4741,I6371);
  not NOT_1176(g6591,I8641);
  not NOT_1177(g5052,I6692);
  not NOT_1178(g6832,I9021);
  not NOT_1179(g4910,I6612);
  not NOT_1180(I2648,g980);
  not NOT_1181(g2234,I3367);
  not NOT_1182(g6853,I9082);
  not NOT_1183(g1890,g1359);
  not NOT_1184(I3883,g2574);
  not NOT_1185(g6420,I8270);
  not NOT_1186(I4240,g2165);
  not NOT_1187(g2330,g1777);
  not NOT_1188(g4108,I5406);
  not NOT_1189(g4609,I6182);
  not NOT_1190(g6507,I8441);
  not NOT_1191(g4308,I5777);
  not NOT_1192(g1011,I2050);
  not NOT_1193(g1734,g952);
  not NOT_1194(I3758,g2041);
  not NOT_1195(g5086,g4732);
  not NOT_1196(g897,g41);
  not NOT_1197(I8040,g6142);
  not NOT_1198(g951,g84);
  not NOT_1199(I8969,g6797);
  not NOT_1200(g2800,g2430);
  not NOT_1201(g5730,I7497);
  not NOT_1202(g2554,I3669);
  not NOT_1203(g4758,I6382);
  not NOT_1204(I2839,g1123);
  not NOT_1205(I3861,g1834);
  not NOT_1206(g6905,I9182);
  not NOT_1207(g3029,I4240);
  not NOT_1208(I3711,g1848);
  not NOT_1209(I9182,g6879);
  not NOT_1210(g3787,I4986);
  not NOT_1211(g2213,I3346);
  not NOT_1212(g5897,g5731);
  not NOT_1213(g5025,g4814);
  not NOT_1214(g6515,g6408);
  not NOT_1215(g4861,I6587);
  not NOT_1216(g5425,I7091);
  not NOT_1217(I4347,g2555);
  not NOT_1218(I2172,g691);
  not NOT_1219(I2278,g917);
  not NOT_1220(g4711,I6315);
  not NOT_1221(g6100,I7796);
  not NOT_1222(I4681,g2947);
  not NOT_1223(g1480,g985);
  not NOT_1224(g2902,g1899);
  not NOT_1225(I8875,g6697);
  not NOT_1226(I2143,g2);
  not NOT_1227(I2343,g1177);
  not NOT_1228(I6139,g4222);
  not NOT_1229(g4133,I5481);
  not NOT_1230(g3297,g3046);
  not NOT_1231(g2512,I3638);
  not NOT_1232(g2090,I3206);
  not NOT_1233(g4846,I6546);
  not NOT_1234(I2134,g705);
  not NOT_1235(I6795,g5022);
  not NOT_1236(I6737,g4662);
  not NOT_1237(I2334,g1193);
  not NOT_1238(I6809,g5051);
  not NOT_1239(I5743,g4022);
  not NOT_1240(g5331,I6995);
  not NOT_1241(I5890,g3878);
  not NOT_1242(I3509,g1461);
  not NOT_1243(g3963,I5217);
  not NOT_1244(g3791,g3388);
  not NOT_1245(I8884,g6704);
  not NOT_1246(I5505,g3860);
  not NOT_1247(g1688,I2688);
  not NOT_1248(I6672,g4752);
  not NOT_1249(g4780,I6434);
  not NOT_1250(g6040,g5824);
  not NOT_1251(g1857,I2961);
  not NOT_1252(I6231,g4350);
  not NOT_1253(I3662,g1688);
  not NOT_1254(g4509,I6039);
  not NOT_1255(g5087,g4736);
  not NOT_1256(I9095,g6855);
  not NOT_1257(g5801,I7600);
  not NOT_1258(g2155,I3274);
  not NOT_1259(I9208,g6922);
  not NOT_1260(g4662,g4640);
  not NOT_1261(I3093,g1426);
  not NOT_1262(g965,I2033);
  not NOT_1263(I3493,g1461);
  not NOT_1264(I3816,g2580);
  not NOT_1265(g1326,g894);
  not NOT_1266(I8235,g6312);
  not NOT_1267(I6099,g4398);
  not NOT_1268(I8282,g6309);
  not NOT_1269(g3049,I4270);
  not NOT_1270(g6528,I8500);
  not NOT_1271(g1760,I2785);
  not NOT_1272(g4493,I6001);
  not NOT_1273(g6351,I8107);
  not NOT_1274(I1850,g210);
  not NOT_1275(g6875,I9092);
  not NOT_1276(g834,g341);
  not NOT_1277(I8988,g6787);
  not NOT_1278(g6530,I8506);
  not NOT_1279(g3575,I4777);
  not NOT_1280(g5045,I6677);
  not NOT_1281(I8693,g6570);
  not NOT_1282(g6655,I8761);
  not NOT_1283(g5445,g5274);
  not NOT_1284(I5713,g4022);
  not NOT_1285(g3604,I4799);
  not NOT_1286(I8548,g6454);
  not NOT_1287(g5491,I7193);
  not NOT_1288(g3498,g2634);
  not NOT_1289(g4381,I5854);
  not NOT_1290(g4847,I6549);
  not NOT_1291(g2118,I3247);
  not NOT_1292(g2619,I3761);
  not NOT_1293(I8555,g6456);
  not NOT_1294(g2367,I3519);
  not NOT_1295(g2872,g1922);
  not NOT_1296(g1608,I2570);
  not NOT_1297(g1220,I2221);
  not NOT_1298(g4700,I6292);
  not NOT_1299(g6410,I8240);
  not NOT_1300(I9164,g6885);
  not NOT_1301(g4397,I5890);
  not NOT_1302(I9233,g6938);
  not NOT_1303(I2776,g1192);
  not NOT_1304(I7640,g5773);
  not NOT_1305(g5407,I7073);
  not NOT_1306(g6884,I9119);
  not NOT_1307(I2593,g1177);
  not NOT_1308(g5059,I6697);
  not NOT_1309(g5920,I7692);
  not NOT_1310(g6839,I9038);
  not NOT_1311(g2457,I3587);
  not NOT_1312(g5578,g5425);
  not NOT_1313(I6444,g4503);
  not NOT_1314(I6269,g4655);
  not NOT_1315(g1423,I2442);
  not NOT_1316(g923,g332);
  not NOT_1317(I5857,g3740);
  not NOT_1318(I7176,g5437);
  not NOT_1319(g1588,g798);
  not NOT_1320(I8113,g6147);
  not NOT_1321(g5582,I7342);
  not NOT_1322(g1161,I2182);
  not NOT_1323(g6278,I7966);
  not NOT_1324(g2686,I3830);
  not NOT_1325(g6372,I8180);
  not NOT_1326(g3162,I4402);
  not NOT_1327(g5261,I6918);
  not NOT_1328(g3019,I4226);
  not NOT_1329(I4294,g2525);
  not NOT_1330(I6543,g4718);
  not NOT_1331(g6618,I8716);
  not NOT_1332(g1665,g985);
  not NOT_1333(I7829,g5926);
  not NOT_1334(I3723,g2158);
  not NOT_1335(g6143,I7865);
  not NOT_1336(g4562,I6132);
  not NOT_1337(g6235,g6062);
  not NOT_1338(g2598,I3726);
  not NOT_1339(g3052,I4273);
  not NOT_1340(g1327,I2334);
  not NOT_1341(I2521,g1063);
  not NOT_1342(I3301,g1730);
  not NOT_1343(g5415,I7081);
  not NOT_1344(g3452,g2625);
  not NOT_1345(g6282,I7996);
  not NOT_1346(I2050,g683);
  not NOT_1347(I5400,g3963);
  not NOT_1348(g6566,I8582);
  not NOT_1349(I8494,g6428);
  not NOT_1350(I4501,g2705);
  not NOT_1351(I6534,g4706);
  not NOT_1352(I8518,g6494);
  not NOT_1353(I3605,g1681);
  not NOT_1354(g4723,I6349);
  not NOT_1355(I8567,g6432);
  not NOT_1356(g4101,I5385);
  not NOT_1357(g6134,I7852);
  not NOT_1358(g5664,g5521);
  not NOT_1359(g2625,I3767);
  not NOT_1360(I7270,g5352);
  not NOT_1361(g2232,I3361);
  not NOT_1362(g6548,I8548);
  not NOT_1363(I6927,g5124);
  not NOT_1364(g3086,I4327);
  not NOT_1365(I2724,g1220);
  not NOT_1366(g2253,I3388);
  not NOT_1367(I2179,g293);
  not NOT_1368(g3486,g2869);
  not NOT_1369(g2813,g2457);
  not NOT_1370(I2379,g1123);
  not NOT_1371(g1696,I2700);
  not NOT_1372(I7073,g5281);
  not NOT_1373(I7796,g5917);
  not NOT_1374(I6885,g4872);
  not NOT_1375(I6414,g4497);
  not NOT_1376(g3504,g2675);
  not NOT_1377(I6946,g5124);
  not NOT_1378(g1732,I2738);
  not NOT_1379(g3881,I5116);
  not NOT_1380(g2740,I3909);
  not NOT_1381(I2658,g1001);
  not NOT_1382(I3441,g1502);
  not NOT_1383(I7069,g5281);
  not NOT_1384(g3070,I4297);
  not NOT_1385(I8264,g6296);
  not NOT_1386(g6621,I8721);
  not NOT_1387(I2835,g1209);
  not NOT_1388(I7469,g5625);
  not NOT_1389(g3897,g3251);
  not NOT_1390(I5023,g3263);
  not NOT_1391(g1472,g952);
  not NOT_1392(g1043,g486);
  not NOT_1393(I5977,g4319);
  not NOT_1394(I8521,g6495);
  not NOT_1395(I6036,g4370);
  not NOT_1396(I8641,g6524);
  not NOT_1397(I2611,g1209);
  not NOT_1398(g893,g23);
  not NOT_1399(g2687,I3833);
  not NOT_1400(I8450,g6412);
  not NOT_1401(I3669,g1739);
  not NOT_1402(g1116,I2154);
  not NOT_1403(g2586,I3711);
  not NOT_1404(I3531,g1593);
  not NOT_1405(I5451,g3967);
  not NOT_1406(I6182,g4249);
  not NOT_1407(g6518,I8470);
  not NOT_1408(g6567,I8585);
  not NOT_1409(I8724,g6533);
  not NOT_1410(I6382,g4460);
  not NOT_1411(g996,I2041);
  not NOT_1412(g3331,g3076);
  not NOT_1413(I3890,g2145);
  not NOT_1414(g4772,I6420);
  not NOT_1415(g5247,g4900);
  not NOT_1416(g4531,I6105);
  not NOT_1417(I5633,g3768);
  not NOT_1418(I8878,g6710);
  not NOT_1419(g1681,I2663);
  not NOT_1420(I3505,g1305);
  not NOT_1421(g6593,I8647);
  not NOT_1422(g3766,I4955);
  not NOT_1423(g1533,g878);
  not NOT_1424(g5564,g5382);
  not NOT_1425(I5103,g3440);
  not NOT_1426(g2525,I3650);
  not NOT_1427(g3801,g3388);
  not NOT_1428(g3487,g2622);
  not NOT_1429(g1914,I3013);
  not NOT_1430(I5696,g3942);
  not NOT_1431(g2691,g2317);
  not NOT_1432(g4011,g3486);
  not NOT_1433(I6798,g5042);
  not NOT_1434(g4856,I6576);
  not NOT_1435(g5741,g5602);
  not NOT_1436(I2802,g1204);
  not NOT_1437(I3074,g1426);
  not NOT_1438(I3474,g1450);
  not NOT_1439(I5753,g4022);
  not NOT_1440(g5638,I7397);
  not NOT_1441(g6160,g5926);
  not NOT_1442(g3226,I4477);
  not NOT_1443(I5508,g3867);
  not NOT_1444(g6360,I8144);
  not NOT_1445(g6933,I9220);
  not NOT_1446(I5944,g4356);
  not NOT_1447(g2962,g2008);
  not NOT_1448(g6521,I8479);
  not NOT_1449(I9098,g6864);
  not NOT_1450(g2158,I3281);
  not NOT_1451(I5472,g3846);
  not NOT_1452(I8981,g6793);
  not NOT_1453(g2506,I3632);
  not NOT_1454(I3080,g1519);
  not NOT_1455(I8674,g6521);
  not NOT_1456(g1820,I2880);
  not NOT_1457(I5043,g3247);
  not NOT_1458(I6495,g4607);
  not NOT_1459(g1936,g1756);
  not NOT_1460(I6437,g4501);
  not NOT_1461(g3173,I4410);
  not NOT_1462(I6102,g4399);
  not NOT_1463(I6302,g4440);
  not NOT_1464(I8997,g6790);
  not NOT_1465(g1117,g32);
  not NOT_1466(I8541,g6452);
  not NOT_1467(g1317,I2306);
  not NOT_1468(g3491,g2608);
  not NOT_1469(g2587,I3714);
  not NOT_1470(I6579,g4798);
  not NOT_1471(I5116,g3259);
  not NOT_1472(I7852,g5993);
  not NOT_1473(I5316,g3557);
  not NOT_1474(g6724,I8866);
  not NOT_1475(I3569,g1789);
  not NOT_1476(g2111,g1384);
  not NOT_1477(g2275,I3422);
  not NOT_1478(g5466,I7146);
  not NOT_1479(I8332,g6306);
  not NOT_1480(g4713,I6321);
  not NOT_1481(I7701,g5720);
  not NOT_1482(g3369,I4646);
  not NOT_1483(I8153,g6185);
  not NOT_1484(g3007,g2197);
  not NOT_1485(g2615,I3755);
  not NOT_1486(g6878,I9101);
  not NOT_1487(I2864,g1177);
  not NOT_1488(g4569,I6143);
  not NOT_1489(g5571,g5395);
  not NOT_1490(g5861,g5636);
  not NOT_1491(g3868,g3491);
  not NOT_1492(g2174,I3313);
  not NOT_1493(g3459,g2664);
  not NOT_1494(g815,I1877);
  not NOT_1495(g1775,g952);
  not NOT_1496(g5448,g5278);
  not NOT_1497(g1922,I3025);
  not NOT_1498(g835,g345);
  not NOT_1499(g5711,I7472);
  not NOT_1500(g6835,I9028);
  not NOT_1501(g1581,g910);
  not NOT_1502(g6882,I9113);
  not NOT_1503(I6042,g4374);
  not NOT_1504(g1060,g107);
  not NOT_1505(g2284,I3431);
  not NOT_1506(I6786,g4824);
  not NOT_1507(g1460,I2457);
  not NOT_1508(g5774,I7517);
  not NOT_1509(g4857,I6579);
  not NOT_1510(g3793,g3491);
  not NOT_1511(g6611,I8699);
  not NOT_1512(g2591,I3720);
  not NOT_1513(g3015,I4220);
  not NOT_1514(g3227,I4480);
  not NOT_1515(g1739,I2749);
  not NOT_1516(I6054,g4194);
  not NOT_1517(g5538,g5331);
  not NOT_1518(I6296,g4436);
  not NOT_1519(I4646,g2602);
  not NOT_1520(I2623,g1161);
  not NOT_1521(g4126,I5460);
  not NOT_1522(g5509,I7251);
  not NOT_1523(g4400,I5899);
  not NOT_1524(g1937,I3044);
  not NOT_1525(g6541,I8535);
  not NOT_1526(I9185,g6877);
  not NOT_1527(I2476,g971);
  not NOT_1528(I7336,g5534);
  not NOT_1529(I8600,g6451);
  not NOT_1530(g2931,g1988);
  not NOT_1531(g4760,I6386);
  not NOT_1532(g1294,I2287);
  not NOT_1533(I1877,g283);
  not NOT_1534(g6332,I8074);
  not NOT_1535(g5067,g4801);
  not NOT_1536(g1190,I2199);
  not NOT_1537(I2175,g25);
  not NOT_1538(g6353,I8113);
  not NOT_1539(g5994,g5873);
  not NOT_1540(I3608,g1461);
  not NOT_1541(g2905,g1994);
  not NOT_1542(I6012,g4167);
  not NOT_1543(g6744,I8910);
  not NOT_1544(I3779,g2125);
  not NOT_1545(g6802,I8972);
  not NOT_1546(g2628,I3770);
  not NOT_1547(g1156,I2175);
  not NOT_1548(g2515,I3641);
  not NOT_1549(g5493,I7197);
  not NOT_1550(I7065,g5281);
  not NOT_1551(g5256,g5077);
  not NOT_1552(I6706,g4731);
  not NOT_1553(g4220,I5644);
  not NOT_1554(g3940,I5177);
  not NOT_1555(I6371,g4569);
  not NOT_1556(I4276,g2170);
  not NOT_1557(g4423,I5920);
  not NOT_1558(I3161,g1270);
  not NOT_1559(I3361,g1331);
  not NOT_1560(g5381,I7039);
  not NOT_1561(g3388,I4667);
  not NOT_1562(I9131,g6855);
  not NOT_1563(I6956,g5124);
  not NOT_1564(g6901,I9170);
  not NOT_1565(I5460,g3771);
  not NOT_1566(I5597,g3821);
  not NOT_1567(I8623,g6542);
  not NOT_1568(g3216,I4459);
  not NOT_1569(I3665,g1824);
  not NOT_1570(g5685,g5552);
  not NOT_1571(g6511,I8453);
  not NOT_1572(I8476,g6457);
  not NOT_1573(I2424,g719);
  not NOT_1574(g743,I1844);
  not NOT_1575(g862,g319);
  not NOT_1576(g2973,I4170);
  not NOT_1577(g1954,I3065);
  not NOT_1578(g3030,I4243);
  not NOT_1579(g1250,g123);
  not NOT_1580(I5739,g3942);
  not NOT_1581(g1363,I2399);
  not NOT_1582(I4986,g3638);
  not NOT_1583(I3999,g1837);
  not NOT_1584(g3247,g2973);
  not NOT_1585(g4127,I5463);
  not NOT_1586(I3346,g1327);
  not NOT_1587(g5950,g5730);
  not NOT_1588(g1053,g197);
  not NOT_1589(g2040,g1738);
  not NOT_1590(g6600,I8668);
  not NOT_1591(g6574,g6484);
  not NOT_1592(I2231,g465);
  not NOT_1593(I1844,g208);
  not NOT_1594(g2440,I3575);
  not NOT_1595(g3564,g2618);
  not NOT_1596(g6714,g6670);
  not NOT_1597(I2643,g965);
  not NOT_1598(g4146,I5520);
  not NOT_1599(I5668,g3828);
  not NOT_1600(g4633,g4284);
  not NOT_1601(I8285,g6310);
  not NOT_1602(I5840,g3732);
  not NOT_1603(I8500,g6431);
  not NOT_1604(g791,I1865);
  not NOT_1605(g4103,I5391);
  not NOT_1606(g6580,g6491);
  not NOT_1607(I7859,g6032);
  not NOT_1608(g5631,g5536);
  not NOT_1609(g3638,g3108);
  not NOT_1610(g5723,I7484);
  not NOT_1611(I9173,g6876);
  not NOT_1612(I3240,g1460);
  not NOT_1613(g4732,I6362);
  not NOT_1614(g3108,I4354);
  not NOT_1615(g3308,g3060);
  not NOT_1616(I6759,g4778);
  not NOT_1617(g2875,g1940);
  not NOT_1618(g4753,I6377);
  not NOT_1619(g4508,I6036);
  not NOT_1620(g917,I1942);
  not NOT_1621(I8809,g6687);
  not NOT_1622(I7342,g5579);
  not NOT_1623(g6623,I8727);
  not NOT_1624(g6076,g5797);
  not NOT_1625(I7081,g5281);
  not NOT_1626(g6889,I9134);
  not NOT_1627(g5751,I7506);
  not NOT_1628(I3316,g1344);
  not NOT_1629(g3589,g3094);
  not NOT_1630(I7481,g5629);
  not NOT_1631(I3034,g1519);
  not NOT_1632(g3466,I4706);
  not NOT_1633(g2410,I3550);
  not NOT_1634(I7692,g5711);
  not NOT_1635(I3434,g1627);
  not NOT_1636(I4516,g2777);
  not NOT_1637(I7497,g5687);
  not NOT_1638(g4116,I5430);
  not NOT_1639(g6375,I8189);
  not NOT_1640(g2884,g1957);
  not NOT_1641(I2044,g681);
  not NOT_1642(g3571,g3084);
  not NOT_1643(g2839,g2535);
  not NOT_1644(g3861,I5084);
  not NOT_1645(g6722,I8860);
  not NOT_1646(g4034,I5333);
  not NOT_1647(I7960,g5925);
  not NOT_1648(g852,g634);
  not NOT_1649(I2269,g899);
  not NOT_1650(g6651,I8749);
  not NOT_1651(g3448,I4684);
  not NOT_1652(g4565,g4195);
  not NOT_1653(I3681,g1821);
  not NOT_1654(I5053,g3710);
  not NOT_1655(g3455,g2637);
  not NOT_1656(g6285,I8005);
  not NOT_1657(g4147,I5523);
  not NOT_1658(g6500,I8420);
  not NOT_1659(g2172,I3307);
  not NOT_1660(I2712,g1203);
  not NOT_1661(I9227,g6937);
  not NOT_1662(I5568,g3897);
  not NOT_1663(g4533,I6111);
  not NOT_1664(g3846,I5053);
  not NOT_1665(g2618,I3758);
  not NOT_1666(I3596,g1305);
  not NOT_1667(g2667,I3811);
  not NOT_1668(g1683,g1017);
  not NOT_1669(g2343,I3493);
  not NOT_1670(g5168,g5099);
  not NOT_1671(I3013,g1519);
  not NOT_1672(g6339,I8093);
  not NOT_1673(g3196,I4433);
  not NOT_1674(g4914,g4816);
  not NOT_1675(g3803,I5002);
  not NOT_1676(g4210,I5630);
  not NOT_1677(I7267,g5458);
  not NOT_1678(g1894,I2989);
  not NOT_1679(I5157,g3454);
  not NOT_1680(g6838,I9035);
  not NOT_1681(I9203,g6921);
  not NOT_1682(I2961,g1731);
  not NOT_1683(g6424,I8282);
  not NOT_1684(g2134,I3258);
  not NOT_1685(I6362,g4569);
  not NOT_1686(g1735,I2745);
  not NOT_1687(I8273,g6301);
  not NOT_1688(g6809,I8981);
  not NOT_1689(g5890,g5753);
  not NOT_1690(g1782,I2828);
  not NOT_1691(I4340,g1935);
  not NOT_1692(I6452,g4629);
  not NOT_1693(I5929,g4152);
  not NOT_1694(g1661,g1076);
  not NOT_1695(I8044,g6252);
  not NOT_1696(g2555,I3672);
  not NOT_1697(g6231,g6044);
  not NOT_1698(g5011,I6649);
  not NOT_1699(I8444,g6421);
  not NOT_1700(g3067,I4294);
  not NOT_1701(I2414,g784);
  not NOT_1702(g729,I1838);
  not NOT_1703(g5411,I7077);
  not NOT_1704(g6523,I8485);
  not NOT_1705(g861,g179);
  not NOT_1706(I2946,g1587);
  not NOT_1707(g2792,g2416);
  not NOT_1708(g1627,I2584);
  not NOT_1709(g4117,I5433);
  not NOT_1710(g1292,I2281);
  not NOT_1711(I5626,g3914);
  not NOT_1712(g3093,I4334);
  not NOT_1713(g898,g47);
  not NOT_1714(g1998,I3109);
  not NOT_1715(g1646,I2617);
  not NOT_1716(g5992,g5869);
  not NOT_1717(g4601,g4191);
  not NOT_1718(g1084,g98);
  not NOT_1719(g6104,I7808);
  not NOT_1720(g854,g646);
  not NOT_1721(g1039,g662);
  not NOT_1722(g1484,I2473);
  not NOT_1723(I3581,g1491);
  not NOT_1724(g6499,I8417);
  not NOT_1725(g1439,I2449);
  not NOT_1726(I9028,g6806);
  not NOT_1727(I8961,g6778);
  not NOT_1728(g4775,I6425);
  not NOT_1729(I6470,g4473);
  not NOT_1730(g5573,g5403);
  not NOT_1731(g3847,I5056);
  not NOT_1732(g5480,I7176);
  not NOT_1733(I6425,g4619);
  not NOT_1734(I2831,g1209);
  not NOT_1735(g2494,I3623);
  not NOT_1736(I2182,g692);
  not NOT_1737(g2518,I3644);
  not NOT_1738(g1583,g1001);
  not NOT_1739(g1702,g1107);
  not NOT_1740(I2382,g719);
  not NOT_1741(I8414,g6418);
  not NOT_1742(g3263,g3015);
  not NOT_1743(I8946,g6778);
  not NOT_1744(g1919,I3022);
  not NOT_1745(I2805,g1205);
  not NOT_1746(I2916,g1643);
  not NOT_1747(g2776,g2378);
  not NOT_1748(I2749,g1209);
  not NOT_1749(g4784,I6444);
  not NOT_1750(g6044,g5824);
  not NOT_1751(g1276,g847);
  not NOT_1752(I4402,g2283);
  not NOT_1753(I3294,g1720);
  not NOT_1754(I3840,g2125);
  not NOT_1755(I6406,g4473);
  not NOT_1756(I5475,g3852);
  not NOT_1757(g6572,I8600);
  not NOT_1758(I4762,g2862);
  not NOT_1759(I7349,g5532);
  not NOT_1760(I6635,g4745);
  not NOT_1761(g2264,I3405);
  not NOT_1762(g6712,g6676);
  not NOT_1763(g851,g606);
  not NOT_1764(I6766,g4783);
  not NOT_1765(I6087,g4392);
  not NOT_1766(I6105,g4400);
  not NOT_1767(g6543,I8541);
  not NOT_1768(g4840,I6528);
  not NOT_1769(I6305,g4441);
  not NOT_1770(I6801,g5045);
  not NOT_1771(g2360,g1793);
  not NOT_1772(g2933,I4123);
  not NOT_1773(g3723,I4903);
  not NOT_1774(g1647,I2620);
  not NOT_1775(g4190,I5600);
  not NOT_1776(I5526,g3848);
  not NOT_1777(I5998,g4157);
  not NOT_1778(I8335,g6308);
  not NOT_1779(I8831,g6665);
  not NOT_1780(I9217,g6931);
  not NOT_1781(g1546,g1101);
  not NOT_1782(I2873,g1161);
  not NOT_1783(I2037,g679);
  not NOT_1784(g6534,I8518);
  not NOT_1785(g6729,I8881);
  not NOT_1786(g3605,I4802);
  not NOT_1787(I5084,g3593);
  not NOT_1788(I5603,g3893);
  not NOT_1789(g2996,I4189);
  not NOT_1790(I2653,g996);
  not NOT_1791(I5484,g3875);
  not NOT_1792(I3942,g1833);
  not NOT_1793(g1503,g878);
  not NOT_1794(I5439,g3730);
  not NOT_1795(I8916,g6742);
  not NOT_1796(g1925,I3028);
  not NOT_1797(I8749,g6560);
  not NOT_1798(g2179,I3328);
  not NOT_1799(g6014,g5824);
  not NOT_1800(g6885,I9122);
  not NOT_1801(I6045,g4375);
  not NOT_1802(g4704,I6302);
  not NOT_1803(g6414,I8252);
  not NOT_1804(I5702,g3845);
  not NOT_1805(g1320,I2315);
  not NOT_1806(g3041,I4258);
  not NOT_1807(g5383,I7045);
  not NOT_1808(g5924,I7704);
  not NOT_1809(g5220,g4903);
  not NOT_1810(I7119,g5303);
  not NOT_1811(g6903,I9176);
  not NOT_1812(g2777,I3965);
  not NOT_1813(g3441,I4681);
  not NOT_1814(g2835,g2506);
  not NOT_1815(I3053,g1407);
  not NOT_1816(I1958,g702);
  not NOT_1817(g4250,I5702);
  not NOT_1818(g6513,I8459);
  not NOT_1819(g913,g658);
  not NOT_1820(I6283,g4613);
  not NOT_1821(I7258,g5458);
  not NOT_1822(I5952,g4367);
  not NOT_1823(g4810,I6488);
  not NOT_1824(g2882,g1854);
  not NOT_1825(I7352,g5533);
  not NOT_1826(g3673,g3075);
  not NOT_1827(I2442,g872);
  not NOT_1828(g1789,I2839);
  not NOT_1829(g6036,g5824);
  not NOT_1830(I8632,g6548);
  not NOT_1831(I2364,g1143);
  not NOT_1832(g980,I2037);
  not NOT_1833(I8653,g6531);
  not NOT_1834(g1771,I2808);
  not NOT_1835(g3772,g3466);
  not NOT_1836(I6582,g4765);
  not NOT_1837(g5051,I6689);
  not NOT_1838(g2981,g2179);
  not NOT_1839(I8579,g6438);
  not NOT_1840(I8869,g6694);
  not NOT_1841(I4489,g2975);
  not NOT_1842(g3458,g2656);
  not NOT_1843(g865,g188);
  not NOT_1844(I2296,g893);
  not NOT_1845(g3890,g3575);
  not NOT_1846(g2997,I4192);
  not NOT_1847(I6015,g4170);
  not NOT_1848(g2541,I3659);
  not NOT_1849(I8752,g6514);
  not NOT_1850(I4471,g3040);
  not NOT_1851(I7170,g5435);
  not NOT_1852(g6422,I8276);
  not NOT_1853(g2353,I3505);
  not NOT_1854(g4929,I6621);
  not NOT_1855(I4955,g3673);
  not NOT_1856(I3626,g1684);
  not NOT_1857(g2744,g2336);
  not NOT_1858(g909,I1935);
  not NOT_1859(g1738,g1108);
  not NOT_1860(g2802,g2437);
  not NOT_1861(g3074,I4303);
  not NOT_1862(g949,g79);
  not NOT_1863(g1991,I3102);
  not NOT_1864(g6560,I8564);
  not NOT_1865(I5320,g3559);
  not NOT_1866(g4626,g4270);
  not NOT_1867(g1340,I2373);
  not NOT_1868(I2029,g677);
  not NOT_1869(I9021,g6812);
  not NOT_1870(g3480,g2986);
  not NOT_1871(g1690,I2692);
  not NOT_1872(g6653,I8755);
  not NOT_1873(g6102,I7802);
  not NOT_1874(I2281,g900);
  not NOT_1875(I7061,g5281);
  not NOT_1876(I7187,g5387);
  not NOT_1877(g6579,g6490);
  not NOT_1878(g5116,g4810);
  not NOT_1879(I5987,g4224);
  not NOT_1880(g5316,I6976);
  not NOT_1881(g1656,I2635);
  not NOT_1882(I6689,g4758);
  not NOT_1883(g5434,I7110);
  not NOT_1884(g2574,I3681);
  not NOT_1885(g2864,g1887);
  not NOT_1886(g4778,I6430);
  not NOT_1887(g855,g650);
  not NOT_1888(g5147,I6809);
  not NOT_1889(I3782,g2145);
  not NOT_1890(g4894,g4813);
  not NOT_1891(I2745,g1249);
  not NOT_1892(I8189,g6179);
  not NOT_1893(I4229,g2284);
  not NOT_1894(I6430,g4620);
  not NOT_1895(g3976,I5252);
  not NOT_1896(I2791,g1236);
  not NOT_1897(I6247,g4609);
  not NOT_1898(I7514,g5590);
  not NOT_1899(I2309,g1236);
  not NOT_1900(I9101,g6855);
  not NOT_1901(g1110,I2140);
  not NOT_1902(I8888,g6708);
  not NOT_1903(g2580,I3691);
  not NOT_1904(g5210,I6874);
  not NOT_1905(g6786,I8946);
  not NOT_1906(I6564,g4712);
  not NOT_1907(I8171,g6170);
  not NOT_1908(I2808,g1161);
  not NOT_1909(I8429,g6425);
  not NOT_1910(g5596,I7358);
  not NOT_1911(g6164,g5926);
  not NOT_1912(g6364,I8156);
  not NOT_1913(g6233,g6052);
  not NOT_1914(I5991,g4226);
  not NOT_1915(I2707,g1190);
  not NOT_1916(g4292,g4059);
  not NOT_1917(I7695,g5714);
  not NOT_1918(I7637,g5751);
  not NOT_1919(g2968,g2179);
  not NOT_1920(I5078,g3719);
  not NOT_1921(g1824,I2890);
  not NOT_1922(g4526,I6090);
  not NOT_1923(I5478,g3859);
  not NOT_1924(g1236,I2234);
  not NOT_1925(I7107,g5277);
  not NOT_1926(I5907,g3883);
  not NOT_1927(g6725,I8869);
  not NOT_1928(g1762,I2791);
  not NOT_1929(g2889,g1975);
  not NOT_1930(I6108,g4403);
  not NOT_1931(g4603,I6170);
  not NOT_1932(g6532,I8512);
  not NOT_1933(I6308,g4443);
  not NOT_1934(I5517,g3885);
  not NOT_1935(I9041,g6835);
  not NOT_1936(I2449,g971);
  not NOT_1937(g4439,I5952);
  not NOT_1938(g5117,I6763);
  not NOT_1939(g6553,I8555);
  not NOT_1940(g4850,I6558);
  not NOT_1941(I8684,g6567);
  not NOT_1942(I5876,g3870);
  not NOT_1943(I8745,g6513);
  not NOT_1944(g2175,I3316);
  not NOT_1945(g2871,g1919);
  not NOT_1946(I2604,g1222);
  not NOT_1947(g3183,I4420);
  not NOT_1948(g2722,I3883);
  not NOT_1949(I4462,g2135);
  not NOT_1950(I8309,g6304);
  not NOT_1951(g1556,g878);
  not NOT_1952(I6066,g4382);
  not NOT_1953(g3779,g3466);
  not NOT_1954(g1222,I2225);
  not NOT_1955(g4702,I6296);
  not NOT_1956(g6412,I8246);
  not NOT_1957(g896,g22);
  not NOT_1958(g3023,g2215);
  not NOT_1959(I7251,g5458);
  not NOT_1960(g1928,I3031);
  not NOT_1961(I7811,g5921);
  not NOT_1962(g6706,I8828);
  not NOT_1963(g5922,I7698);
  not NOT_1964(I8707,g6520);
  not NOT_1965(g1064,g102);
  not NOT_1966(I2584,g839);
  not NOT_1967(I5214,g3567);
  not NOT_1968(g6888,I9131);
  not NOT_1969(g1899,I2998);
  not NOT_1970(I6048,g4376);
  not NOT_1971(g5581,I7339);
  not NOT_1972(I6448,g4626);
  not NOT_1973(g6371,I8177);
  not NOT_1974(g4276,I5731);
  not NOT_1975(I4249,g2525);
  not NOT_1976(g5597,I7361);
  not NOT_1977(I3004,g1426);
  not NOT_1978(I1825,g361);
  not NOT_1979(g4561,g4189);
  not NOT_1980(g2838,g2515);
  not NOT_1981(I3647,g1747);
  not NOT_1982(g3451,g2615);
  not NOT_1983(I2162,g197);
  not NOT_1984(g1563,g1006);
  not NOT_1985(I9011,g6819);
  not NOT_1986(I4192,g1847);
  not NOT_1987(g2809,I4019);
  not NOT_1988(I3764,g2044);
  not NOT_1989(g5784,I7583);
  not NOT_1990(I3546,g1586);
  not NOT_1991(I5002,g3612);
  not NOT_1992(g4527,I6093);
  not NOT_1993(g4404,I5907);
  not NOT_1994(g1295,I2290);
  not NOT_1995(g4647,g4296);
  not NOT_1996(g3346,I4623);
  not NOT_1997(I5236,g3545);
  not NOT_1998(g2672,I3816);
  not NOT_1999(g2231,I3358);
  not NOT_2000(g4764,I6400);
  not NOT_2001(g5995,g5824);
  not NOT_2002(I9074,g6844);
  not NOT_2003(g5479,I7173);
  not NOT_2004(g2643,I3785);
  not NOT_2005(I6780,g4825);
  not NOT_2006(g6745,I8913);
  not NOT_2007(g1394,g1206);
  not NOT_2008(g4503,I6023);
  not NOT_2009(I7612,g5605);
  not NOT_2010(g1731,I2735);
  not NOT_2011(I2728,g1232);
  not NOT_2012(g1557,g1017);
  not NOT_2013(g2634,I3776);
  not NOT_2014(g1966,I3077);
  not NOT_2015(g4224,g4046);
  not NOT_2016(I5556,g4059);
  not NOT_2017(I2185,g29);
  not NOT_2018(g2104,g1372);
  not NOT_2019(g2099,g1366);
  not NOT_2020(g3240,I4519);
  not NOT_2021(I2385,g784);
  not NOT_2022(g6707,I8831);
  not NOT_2023(g1471,I2464);
  not NOT_2024(g4120,I5442);
  not NOT_2025(I4031,g1846);
  not NOT_2026(g4320,g4011);
  not NOT_2027(I4252,g2555);
  not NOT_2028(I3617,g1305);
  not NOT_2029(I3906,g2234);
  not NOT_2030(I6093,g4394);
  not NOT_2031(I8162,g6189);
  not NOT_2032(g3043,I4264);
  not NOT_2033(g971,g658);
  not NOT_2034(I5899,g3748);
  not NOT_2035(I4176,g2268);
  not NOT_2036(I6816,g5111);
  not NOT_2037(I3516,g1295);
  not NOT_2038(g2754,g2347);
  not NOT_2039(g4617,g4242);
  not NOT_2040(g3034,I4249);
  not NOT_2041(g1254,g152);
  not NOT_2042(g1814,I2873);
  not NOT_2043(g6575,g6486);
  not NOT_2044(g4516,I6060);
  not NOT_2045(g6715,g6673);
  not NOT_2046(g4771,I6417);
  not NOT_2047(g2044,I3161);
  not NOT_2048(I6685,g4716);
  not NOT_2049(g5250,g4929);
  not NOT_2050(g6604,I8678);
  not NOT_2051(g1038,g127);
  not NOT_2052(I6397,g4473);
  not NOT_2053(g6498,I8414);
  not NOT_2054(g1773,I2814);
  not NOT_2055(I2131,g24);
  not NOT_2056(g5432,I7104);
  not NOT_2057(g4299,I5756);
  not NOT_2058(g6833,I9024);
  not NOT_2059(I8730,g6535);
  not NOT_2060(g5453,g5296);
  not NOT_2061(I4270,g2555);
  not NOT_2062(g2862,I4066);
  not NOT_2063(I2635,g1055);
  not NOT_2064(g2712,g2320);
  not NOT_2065(I8881,g6711);
  not NOT_2066(I5394,g4016);
  not NOT_2067(g1769,I2802);
  not NOT_2068(g3914,I5153);
  not NOT_2069(g6584,I8620);
  not NOT_2070(I1859,g277);
  not NOT_2071(g6539,I8531);
  not NOT_2072(g6896,I9155);
  not NOT_2073(g1836,I2922);
  not NOT_2074(g5568,g5423);
  not NOT_2075(I8070,g6116);
  not NOT_2076(I5731,g3942);
  not NOT_2077(I8470,g6461);
  not NOT_2078(I8897,g6707);
  not NOT_2079(g1918,I3019);
  not NOT_2080(I3244,g1772);
  not NOT_2081(I7490,g5583);
  not NOT_2082(I4980,g3546);
  not NOT_2083(g5912,g5853);
  not NOT_2084(I4324,g1918);
  not NOT_2085(I3140,g1317);
  not NOT_2086(g2961,g1861);
  not NOT_2087(I5071,g3263);
  not NOT_2088(I3340,g1282);
  not NOT_2089(I5705,g3942);
  not NOT_2090(g6162,g5926);
  not NOT_2091(I3478,g1450);
  not NOT_2092(g6362,I8150);
  not NOT_2093(g6419,I8267);
  not NOT_2094(I6723,g4761);
  not NOT_2095(g4140,I5502);
  not NOT_2096(g6052,g5824);
  not NOT_2097(g2927,g1979);
  not NOT_2098(I5948,g4360);
  not NOT_2099(I9220,g6930);
  not NOT_2100(g2885,g1963);
  not NOT_2101(I7355,g5535);
  not NOT_2102(I8678,g6565);
  not NOT_2103(I2445,g971);
  not NOT_2104(g2660,I3804);
  not NOT_2105(g2946,g2296);
  not NOT_2106(g938,g59);
  not NOT_2107(g4435,I5944);
  not NOT_2108(I2373,g1143);
  not NOT_2109(g4517,I6063);
  not NOT_2110(I7698,g5717);
  not NOT_2111(I3656,g1484);
  not NOT_2112(g3601,I4794);
  not NOT_2113(I2491,g821);
  not NOT_2114(g2903,g1902);
  not NOT_2115(I8635,g6552);
  not NOT_2116(g6728,I8878);
  not NOT_2117(g6486,g6363);
  not NOT_2118(I2169,g269);
  not NOT_2119(g942,g69);
  not NOT_2120(g6730,I8884);
  not NOT_2121(I9161,g6880);
  not NOT_2122(g3775,g3388);
  not NOT_2123(g6504,I8432);
  not NOT_2124(g3922,I5157);
  not NOT_2125(I7463,g5622);
  not NOT_2126(I2578,g1209);
  not NOT_2127(g6385,g6271);
  not NOT_2128(g6881,I9110);
  not NOT_2129(I5409,g3980);
  not NOT_2130(g2036,g1764);
  not NOT_2131(g706,I1825);
  not NOT_2132(I6441,g4624);
  not NOT_2133(g4915,g4669);
  not NOT_2134(g2178,I3325);
  not NOT_2135(g2436,I3569);
  not NOT_2136(g2679,I3823);
  not NOT_2137(g6070,g5824);
  not NOT_2138(g2378,I3525);
  not NOT_2139(g3060,I4285);
  not NOT_2140(I3310,g1640);
  not NOT_2141(g6897,I9158);
  not NOT_2142(g1837,I2925);
  not NOT_2143(I8755,g6561);
  not NOT_2144(g3460,g2667);
  not NOT_2145(I8226,g6328);
  not NOT_2146(g6425,I8285);
  not NOT_2147(g2135,I3261);
  not NOT_2148(I4510,g2753);
  not NOT_2149(I9146,g6890);
  not NOT_2150(g4110,I5412);
  not NOT_2151(I7167,g5434);
  not NOT_2152(I7318,g5452);
  not NOT_2153(I4291,g2241);
  not NOT_2154(g5894,g5731);
  not NOT_2155(g2805,g2443);
  not NOT_2156(g910,I1938);
  not NOT_2157(g1788,g985);
  not NOT_2158(g2422,I3560);
  not NOT_2159(I6772,g4788);
  not NOT_2160(I7193,g5466);
  not NOT_2161(I8491,g6480);
  not NOT_2162(g3079,I4312);
  not NOT_2163(I6531,g4704);
  not NOT_2164(g4402,g4017);
  not NOT_2165(g784,I1862);
  not NOT_2166(g1249,I2240);
  not NOT_2167(g4824,g4615);
  not NOT_2168(g837,g353);
  not NOT_2169(g5661,g5518);
  not NOT_2170(g3840,I5043);
  not NOT_2171(g719,I1835);
  not NOT_2172(I3590,g1781);
  not NOT_2173(g6406,I8232);
  not NOT_2174(g5475,I7161);
  not NOT_2175(I7686,g5705);
  not NOT_2176(g1842,g1612);
  not NOT_2177(I2721,g1219);
  not NOT_2178(g1192,g44);
  not NOT_2179(I8459,g6427);
  not NOT_2180(g6105,I7811);
  not NOT_2181(g6087,g5813);
  not NOT_2182(g6801,I8969);
  not NOT_2183(g6305,I8027);
  not NOT_2184(g5292,I6942);
  not NOT_2185(I8767,g6619);
  not NOT_2186(g6487,g6365);
  not NOT_2187(I3556,g1484);
  not NOT_2188(g3501,g2650);
  not NOT_2189(I3222,g1790);
  not NOT_2190(I8535,g6447);
  not NOT_2191(g4657,I6244);
  not NOT_2192(I8582,g6439);
  not NOT_2193(g1854,I2958);
  not NOT_2194(I9116,g6864);
  not NOT_2195(I8261,g6298);
  not NOT_2196(g5084,g4727);
  not NOT_2197(g4222,I5654);
  not NOT_2198(g2437,I3572);
  not NOT_2199(g2653,I3797);
  not NOT_2200(I6992,g5151);
  not NOT_2201(I1932,g667);
  not NOT_2202(g2102,I3222);
  not NOT_2203(g5439,g5261);
  not NOT_2204(I3785,g2346);
  not NOT_2205(I2940,g1653);
  not NOT_2206(I5837,g3850);
  not NOT_2207(g2869,g2433);
  not NOT_2208(I2388,g878);
  not NOT_2209(I6573,g4721);
  not NOT_2210(I3563,g1461);
  not NOT_2211(g5702,I7463);
  not NOT_2212(I8246,g6290);
  not NOT_2213(g1219,I2218);
  not NOT_2214(g1640,I2601);
  not NOT_2215(g2752,g2343);
  not NOT_2216(g6373,I8183);
  not NOT_2217(g3363,g3110);
  not NOT_2218(g6491,g6373);
  not NOT_2219(g5919,I7689);
  not NOT_2220(I2671,g1017);
  not NOT_2221(g1812,I2867);
  not NOT_2222(I8721,g6534);
  not NOT_2223(I2428,g774);
  not NOT_2224(g4563,g4190);
  not NOT_2225(g3053,I4276);
  not NOT_2226(g1176,I2190);
  not NOT_2227(g2265,I3408);
  not NOT_2228(g3453,g2628);
  not NOT_2229(g6283,I7999);
  not NOT_2230(g6369,I8171);
  not NOT_2231(g2042,I3155);
  not NOT_2232(g6602,I8674);
  not NOT_2233(I5249,g3589);
  not NOT_2234(g6407,I8235);
  not NOT_2235(g6578,g6489);
  not NOT_2236(g4844,I6540);
  not NOT_2237(g2164,I3291);
  not NOT_2238(g1286,g854);
  not NOT_2239(g2364,I3516);
  not NOT_2240(g2233,I3364);
  not NOT_2241(g4194,I5612);
  not NOT_2242(g1911,I3010);
  not NOT_2243(g4394,I5885);
  not NOT_2244(g6535,I8521);
  not NOT_2245(I6976,g5136);
  not NOT_2246(g3912,g3505);
  not NOT_2247(I2741,g1222);
  not NOT_2248(g5527,I7267);
  not NOT_2249(g6582,I8614);
  not NOT_2250(I8940,g6783);
  not NOT_2251(g4731,I6359);
  not NOT_2252(I2910,g1645);
  not NOT_2253(I3071,g1504);
  not NOT_2254(g5647,g5509);
  not NOT_2255(I3705,g2316);
  not NOT_2256(I3471,g1450);
  not NOT_2257(g2296,I3441);
  not NOT_2258(g1733,I2741);
  not NOT_2259(I2638,g1123);
  not NOT_2260(g1270,g844);
  not NOT_2261(g5546,g5388);
  not NOT_2262(I5854,g3857);
  not NOT_2263(I4465,g2945);
  not NOT_2264(g6015,g5857);
  not NOT_2265(g4705,I6305);
  not NOT_2266(g6415,I8255);
  not NOT_2267(I6126,g4240);
  not NOT_2268(I6400,g4473);
  not NOT_2269(g4242,I5686);
  not NOT_2270(I2883,g1143);
  not NOT_2271(I8671,g6519);
  not NOT_2272(g5925,I7707);
  not NOT_2273(I8030,g6239);
  not NOT_2274(I4433,g2103);
  not NOT_2275(g1324,I2327);
  not NOT_2276(I5708,g3942);
  not NOT_2277(I5520,g3835);
  not NOT_2278(g6721,I8857);
  not NOT_2279(I5640,g3770);
  not NOT_2280(g5120,I6772);
  not NOT_2281(I8564,g6429);
  not NOT_2282(g2706,I3861);
  not NOT_2283(I5252,g3546);
  not NOT_2284(I3773,g2524);
  not NOT_2285(g1177,I2193);
  not NOT_2286(g4150,I5532);
  not NOT_2287(I2165,g690);
  not NOT_2288(g1206,I2212);
  not NOT_2289(g4350,g4010);
  not NOT_2290(g2888,g1972);
  not NOT_2291(I7358,g5565);
  not NOT_2292(I4195,g2173);
  not NOT_2293(g2029,I3134);
  not NOT_2294(I7506,g5584);
  not NOT_2295(I5376,g4014);
  not NOT_2296(g2171,I3304);
  not NOT_2297(I4337,g1934);
  not NOT_2298(I8910,g6730);
  not NOT_2299(g2787,g2405);
  not NOT_2300(g6502,I8426);
  not NOT_2301(g2956,g1861);
  not NOT_2302(I6023,g4151);
  not NOT_2303(I8638,g6553);
  not NOT_2304(g1287,g855);
  not NOT_2305(g2675,I3819);
  not NOT_2306(I3836,g1832);
  not NOT_2307(I3212,g1806);
  not NOT_2308(I7587,g5605);
  not NOT_2309(g6940,I9233);
  not NOT_2310(g4769,g4606);
  not NOT_2311(g1849,I2949);
  not NOT_2312(g3778,g3388);
  not NOT_2313(g6188,g5950);
  not NOT_2314(I2196,g3);
  not NOT_2315(g5299,I6949);
  not NOT_2316(g1781,I2825);
  not NOT_2317(I6051,g4185);
  not NOT_2318(g1898,I2995);
  not NOT_2319(g3782,g3388);
  not NOT_2320(I8217,g6319);
  not NOT_2321(I8758,g6562);
  not NOT_2322(I8066,g6114);
  not NOT_2323(g5892,g5742);
  not NOT_2324(I6327,g4451);
  not NOT_2325(g6428,I8290);
  not NOT_2326(g3075,I4306);
  not NOT_2327(g4229,g4059);
  not NOT_2328(g2109,I3235);
  not NOT_2329(I7284,g5383);
  not NOT_2330(I4255,g2179);
  not NOT_2331(I6346,g4563);
  not NOT_2332(I8165,g6189);
  not NOT_2333(g4822,g4614);
  not NOT_2334(g1291,I2278);
  not NOT_2335(I5124,g3719);
  not NOT_2336(I2067,g686);
  not NOT_2337(g6564,I8576);
  not NOT_2338(I5324,g3466);
  not NOT_2339(I7832,g5943);
  not NOT_2340(g6826,I9011);
  not NOT_2341(I5469,g3838);
  not NOT_2342(I2290,g971);
  not NOT_2343(g1344,I2379);
  not NOT_2344(I4354,g1953);
  not NOT_2345(g5140,I6798);
  not NOT_2346(I5177,g3267);
  not NOT_2347(g3084,I4321);
  not NOT_2348(g5478,I7170);
  not NOT_2349(g1819,I2877);
  not NOT_2350(I6753,g4772);
  not NOT_2351(g2957,g1861);
  not NOT_2352(I8803,g6685);
  not NOT_2353(g1088,I2119);
  not NOT_2354(g1852,I2952);
  not NOT_2355(I6072,g4385);
  not NOT_2356(g6609,I8693);
  not NOT_2357(g5435,I7113);
  not NOT_2358(g6308,I8034);
  not NOT_2359(I3062,g1776);
  not NOT_2360(g5082,g4723);
  not NOT_2361(g2449,I3584);
  not NOT_2362(I3620,g1484);
  not NOT_2363(I3462,g1450);
  not NOT_2364(I8538,g6450);
  not NOT_2365(g2575,I3684);
  not NOT_2366(g2865,g2296);
  not NOT_2367(g6883,I9116);
  not NOT_2368(g5876,I7640);
  not NOT_2369(g4837,g4473);
  not NOT_2370(I8509,g6437);
  not NOT_2371(I2700,g1173);
  not NOT_2372(g2604,I3736);
  not NOT_2373(I4267,g2525);
  not NOT_2374(g2098,g1363);
  not NOT_2375(I4312,g2555);
  not NOT_2376(g4620,g4251);
  not NOT_2377(g4462,I5977);
  not NOT_2378(g6589,I8635);
  not NOT_2379(g945,g536);
  not NOT_2380(I8662,g6525);
  not NOT_2381(I3788,g2554);
  not NOT_2382(g6466,I8332);
  not NOT_2383(g5915,I7679);
  not NOT_2384(g3952,I5182);
  not NOT_2385(I6434,g4622);
  not NOT_2386(I8467,g6457);
  not NOT_2387(I8994,g6789);
  not NOT_2388(I8290,g6291);
  not NOT_2389(g1114,I2150);
  not NOT_2390(g6165,g5926);
  not NOT_2391(g6571,I8597);
  not NOT_2392(g6365,I8159);
  not NOT_2393(g2584,I3705);
  not NOT_2394(g4788,I6452);
  not NOT_2395(g6048,g5824);
  not NOT_2396(I1841,g207);
  not NOT_2397(g6711,I8843);
  not NOT_2398(I8093,g6122);
  not NOT_2399(g5110,I6740);
  not NOT_2400(g4249,I5699);
  not NOT_2401(g5310,g5067);
  not NOT_2402(I3298,g1725);
  not NOT_2403(g1825,I2893);
  not NOT_2404(g6827,I9014);
  not NOT_2405(g1650,I2627);
  not NOT_2406(I3485,g1450);
  not NOT_2407(g3527,I4743);
  not NOT_2408(g809,I1874);
  not NOT_2409(I6697,g4722);
  not NOT_2410(g4842,I6534);
  not NOT_2411(g849,g598);
  not NOT_2412(g2268,I3419);
  not NOT_2413(g4192,I5606);
  not NOT_2414(g4392,I5879);
  not NOT_2415(g3546,g3095);
  not NOT_2416(g4485,I5987);
  not NOT_2417(I2817,g1222);
  not NOT_2418(g5824,g5631);
  not NOT_2419(g1336,I2361);
  not NOT_2420(g6803,I8975);
  not NOT_2421(g3970,I5236);
  not NOT_2422(g1594,g1143);
  not NOT_2423(g4854,I6570);
  not NOT_2424(g6538,g6469);
  not NOT_2425(g1972,I3083);
  not NOT_2426(I5923,g4299);
  not NOT_2427(g6509,I8447);
  not NOT_2428(g1806,I2857);
  not NOT_2429(g5877,I7643);
  not NOT_2430(g5590,I7352);
  not NOT_2431(g1943,I3050);
  not NOT_2432(I3708,g1946);
  not NOT_2433(g3224,I4471);
  not NOT_2434(g2086,I3198);
  not NOT_2435(g2728,I3890);
  not NOT_2436(I3031,g1504);
  not NOT_2437(I4468,g2583);
  not NOT_2438(g3320,g3067);
  not NOT_2439(g6067,g5788);
  not NOT_2440(g1887,I2982);
  not NOT_2441(I3431,g1275);
  not NOT_2442(g1122,I2162);
  not NOT_2443(g6418,I8264);
  not NOT_2444(g6467,I8335);
  not NOT_2445(g1322,I2321);
  not NOT_2446(g4520,I6072);
  not NOT_2447(g1934,I3037);
  not NOT_2448(I2041,g680);
  not NOT_2449(I3376,g1328);
  not NOT_2450(g4431,I5938);
  not NOT_2451(g4252,I5708);
  not NOT_2452(I1874,g282);
  not NOT_2453(I3405,g1321);
  not NOT_2454(g3906,g3575);
  not NOT_2455(g2470,I3602);
  not NOT_2456(g3789,g3388);
  not NOT_2457(g5064,I6706);
  not NOT_2458(g2025,g1276);
  not NOT_2459(g6493,g6375);
  not NOT_2460(g5899,g5753);
  not NOT_2461(I6775,g4790);
  not NOT_2462(g4376,I5843);
  not NOT_2463(g4405,I5910);
  not NOT_2464(g3771,I4964);
  not NOT_2465(I5825,g3914);
  not NOT_2466(g872,g143);
  not NOT_2467(g1550,g996);
  not NOT_2468(I6060,g4380);
  not NOT_2469(g4286,I5743);
  not NOT_2470(g4765,I6403);
  not NOT_2471(I1880,g276);
  not NOT_2472(I4198,g2276);
  not NOT_2473(g3299,g3049);
  not NOT_2474(g5563,g5381);
  not NOT_2475(I4398,g2086);
  not NOT_2476(g4911,I6615);
  not NOT_2477(I3733,g2031);
  not NOT_2478(g6700,I8818);
  not NOT_2479(g1395,I2428);
  not NOT_2480(g1891,I2986);
  not NOT_2481(g1337,I2364);
  not NOT_2482(g5237,g5083);
  not NOT_2483(g3892,g3575);
  not NOT_2484(g2678,g2312);
  not NOT_2485(I3225,g1813);
  not NOT_2486(g6421,I8273);
  not NOT_2487(I2890,g1123);
  not NOT_2488(I8585,g6442);
  not NOT_2489(I5594,g3821);
  not NOT_2490(g4270,I5723);
  not NOT_2491(I7372,g5493);
  not NOT_2492(g1807,I2860);
  not NOT_2493(g4225,g4059);
  not NOT_2494(g2682,I3826);
  not NOT_2495(g2766,g2361);
  not NOT_2496(I6995,g5220);
  not NOT_2497(I1935,g666);
  not NOT_2498(g2087,g1352);
  not NOT_2499(g2105,g1375);
  not NOT_2500(I6937,g5124);
  not NOT_2501(I7143,g5323);
  not NOT_2502(I8441,g6419);
  not NOT_2503(g2801,I4003);
  not NOT_2504(I2411,g736);
  not NOT_2505(g5089,I6723);
  not NOT_2506(g5489,I7187);
  not NOT_2507(I5065,g3714);
  not NOT_2508(g4124,I5454);
  not NOT_2509(g714,g131);
  not NOT_2510(I3540,g1670);
  not NOT_2511(g4980,g4678);
  not NOT_2512(g2748,I3923);
  not NOT_2513(g6562,I8570);
  not NOT_2514(I3206,g1823);
  not NOT_2515(g5705,I7466);
  not NOT_2516(I2992,g1741);
  not NOT_2517(g3478,g2695);
  not NOT_2518(g1142,I2169);
  not NOT_2519(g2755,g2350);
  not NOT_2520(I4258,g2169);
  not NOT_2521(g5242,g5085);
  not NOT_2522(I8168,g6170);
  not NOT_2523(g6723,I8863);
  not NOT_2524(g1255,g161);
  not NOT_2525(I5033,g3527);
  not NOT_2526(g6101,I7799);
  not NOT_2527(g6817,I8988);
  not NOT_2528(I5433,g3728);
  not NOT_2529(g4206,I5626);
  not NOT_2530(g3082,I4315);
  not NOT_2531(g3482,g2713);
  not NOT_2532(I8531,g6444);
  not NOT_2533(g1692,I2696);
  not NOT_2534(g6605,I8681);
  not NOT_2535(g1726,I2728);
  not NOT_2536(g3876,I5109);
  not NOT_2537(g2173,I3310);
  not NOT_2538(I6942,g5124);
  not NOT_2539(g2091,g1355);
  not NOT_2540(I5496,g3839);
  not NOT_2541(g1960,I3071);
  not NOT_2542(g2491,I3620);
  not NOT_2543(g5150,I6816);
  not NOT_2544(g4849,I6555);
  not NOT_2545(g2169,I3298);
  not NOT_2546(g2283,I3428);
  not NOT_2547(I7113,g5295);
  not NOT_2548(I8411,g6415);
  not NOT_2549(I5337,g3564);
  not NOT_2550(I5913,g3751);
  not NOT_2551(g2602,g2061);
  not NOT_2552(g6585,I8623);
  not NOT_2553(g2007,g1411);
  not NOT_2554(g5773,I7514);
  not NOT_2555(g4399,I5896);
  not NOT_2556(I3797,g2125);
  not NOT_2557(I6250,g4514);
  not NOT_2558(g2059,g1402);
  not NOT_2559(g2920,g1947);
  not NOT_2560(I4170,g2157);
  not NOT_2561(g4781,I6437);
  not NOT_2562(g6441,I8309);
  not NOT_2563(I8074,g6118);
  not NOT_2564(g2767,g2364);
  not NOT_2565(g4900,I6607);
  not NOT_2566(g1783,I2831);
  not NOT_2567(g3110,I4358);
  not NOT_2568(I4821,g2877);
  not NOT_2569(I2688,g1030);
  not NOT_2570(I2857,g1161);
  not NOT_2571(g2535,I3653);
  not NOT_2572(I3291,g1714);
  not NOT_2573(g1979,I3090);
  not NOT_2574(g1112,g336);
  not NOT_2575(g1267,g843);
  not NOT_2576(I7494,g5691);
  not NOT_2577(g4510,I6042);
  not NOT_2578(I3144,g1319);
  not NOT_2579(g5918,I7686);
  not NOT_2580(g1001,I2044);
  not NOT_2581(g3002,g2215);
  not NOT_2582(I8573,g6435);
  not NOT_2583(I8863,g6700);
  not NOT_2584(I4483,g3082);
  not NOT_2585(g1293,I2284);
  not NOT_2586(g6368,I8168);
  not NOT_2587(g4144,I5514);
  not NOT_2588(I8713,g6522);
  not NOT_2589(I7593,g5605);
  not NOT_2590(I3819,g2044);
  not NOT_2591(g3236,I4507);
  not NOT_2592(g1329,I2340);
  not NOT_2593(I3694,g1811);
  not NOT_2594(g1761,I2788);
  not NOT_2595(g857,g170);
  not NOT_2596(g5993,g5872);
  not NOT_2597(g6531,I8509);
  not NOT_2598(I5081,g3589);
  not NOT_2599(I3923,g2581);
  not NOT_2600(I4306,g1898);
  not NOT_2601(I2760,g1193);
  not NOT_2602(g2664,I3808);
  not NOT_2603(I5481,g3866);
  not NOT_2604(I3488,g1295);
  not NOT_2605(g6743,I8907);
  not NOT_2606(g6890,I9137);
  not NOT_2607(g1830,I2904);
  not NOT_2608(I5692,g3942);
  not NOT_2609(I7264,g5458);
  not NOT_2610(g4852,I6564);
  not NOT_2611(g6505,I8435);
  not NOT_2612(I3215,g1820);
  not NOT_2613(g1221,g46);
  not NOT_2614(g6411,I8243);
  not NOT_2615(g6734,I8894);
  not NOT_2616(g3222,I4465);
  not NOT_2617(I3886,g2215);
  not NOT_2618(I8857,g6698);
  not NOT_2619(g1703,I2707);
  not NOT_2620(I2608,g1143);
  not NOT_2621(g5921,I7695);
  not NOT_2622(g4215,I5637);
  not NOT_2623(I2779,g1038);
  not NOT_2624(I7996,g6137);
  not NOT_2625(g6074,g5794);
  not NOT_2626(g3064,I4291);
  not NOT_2627(g3785,g3466);
  not NOT_2628(g1624,I2581);
  not NOT_2629(g1953,I3062);
  not NOT_2630(I4003,g2284);
  not NOT_2631(g5895,g5742);
  not NOT_2632(g4114,I5424);
  not NOT_2633(g4314,g4080);
  not NOT_2634(I2588,g1193);
  not NOT_2635(I3650,g1650);
  not NOT_2636(g6080,g5805);
  not NOT_2637(I2361,g1075);
  not NOT_2638(g6573,I8603);
  not NOT_2639(I4391,g2275);
  not NOT_2640(g6713,g6679);
  not NOT_2641(I3408,g1644);
  not NOT_2642(g3237,I4510);
  not NOT_2643(I7835,g5926);
  not NOT_2644(I2327,g1222);
  not NOT_2645(g6569,I8591);
  not NOT_2646(g2030,I3137);
  not NOT_2647(g5788,I7587);
  not NOT_2648(g2430,I3563);
  not NOT_2649(I2346,g1193);
  not NOT_2650(g4136,I5490);
  not NOT_2651(I8183,g6176);
  not NOT_2652(I4223,g2176);
  not NOT_2653(I8220,g6322);
  not NOT_2654(g4768,I6410);
  not NOT_2655(g1848,I2946);
  not NOT_2656(I9140,g6888);
  not NOT_2657(g2826,g2481);
  not NOT_2658(g1699,I2703);
  not NOT_2659(g1747,I2760);
  not NOT_2660(g838,g564);
  not NOT_2661(I6075,g4386);
  not NOT_2662(I2696,g1156);
  not NOT_2663(I4757,g2861);
  not NOT_2664(I7799,g5918);
  not NOT_2665(I3065,g1426);
  not NOT_2666(g3557,g2598);
  not NOT_2667(I5746,g4022);
  not NOT_2668(g4806,g4473);
  not NOT_2669(g5392,I7058);
  not NOT_2670(I8423,g6423);
  not NOT_2671(I9035,g6812);
  not NOT_2672(I6949,g5050);
  not NOT_2673(g4943,I6635);
  not NOT_2674(I3465,g1724);
  not NOT_2675(I3322,g1333);
  not NOT_2676(I9082,g6849);
  not NOT_2677(g3705,g3014);
  not NOT_2678(I8588,g6443);
  not NOT_2679(I4522,g2801);
  not NOT_2680(I2753,g1174);
  not NOT_2681(g842,g571);
  not NOT_2682(I6292,g4434);
  not NOT_2683(I4315,g2245);
  not NOT_2684(g3242,g3083);
  not NOT_2685(g4122,I5448);
  not NOT_2686(g4228,I5668);
  not NOT_2687(g4322,I5793);
  not NOT_2688(I2240,g19);
  not NOT_2689(I1938,g332);
  not NOT_2690(g2108,I3232);
  not NOT_2691(g2609,I3749);
  not NOT_2692(I6646,g4687);
  not NOT_2693(g2308,I3452);
  not NOT_2694(I8665,g6527);
  not NOT_2695(I8051,g6108);
  not NOT_2696(I7153,g5358);
  not NOT_2697(g2883,g1954);
  not NOT_2698(I6084,g4391);
  not NOT_2699(I6039,g4182);
  not NOT_2700(I5068,g3571);
  not NOT_2701(I3096,g1439);
  not NOT_2702(g1644,I2611);
  not NOT_2703(I3496,g1326);
  not NOT_2704(g715,g135);
  not NOT_2705(I3550,g1295);
  not NOT_2706(I7802,g5920);
  not NOT_2707(g5708,I7469);
  not NOT_2708(g1119,I2159);
  not NOT_2709(g1319,I2312);
  not NOT_2710(g2066,g1341);
  not NOT_2711(g3150,I4391);
  not NOT_2712(g5219,I6885);
  not NOT_2713(I3137,g1315);
  not NOT_2714(I8103,g6134);
  not NOT_2715(I3395,g1286);
  not NOT_2716(I3337,g1338);
  not NOT_2717(g4496,I6008);
  not NOT_2718(g1352,I2391);
  not NOT_2719(I9110,g6864);
  not NOT_2720(g1577,g1001);
  not NOT_2721(g4550,I6126);
  not NOT_2722(g3773,g3466);
  not NOT_2723(g4845,I6543);
  not NOT_2724(I4537,g2877);
  not NOT_2725(I8696,g6569);
  not NOT_2726(g2165,I3294);
  not NOT_2727(g5958,g5818);
  not NOT_2728(I2147,g6);
  not NOT_2729(g6608,I8690);
  not NOT_2730(g4195,I5615);
  not NOT_2731(g4137,I5493);
  not NOT_2732(g830,g338);
  not NOT_2733(I5716,g3942);
  not NOT_2734(g3769,g3622);
  not NOT_2735(I9002,g6802);
  not NOT_2736(g2827,g2485);
  not NOT_2737(I6952,g5124);
  not NOT_2738(I5848,g3856);
  not NOT_2739(g3836,I5033);
  not NOT_2740(g3212,I4455);
  not NOT_2741(g6423,I8279);
  not NOT_2742(I4243,g1853);
  not NOT_2743(g2333,I3485);
  not NOT_2744(I8240,g6287);
  not NOT_2745(g1975,I3086);
  not NOT_2746(I5699,g3844);
  not NOT_2747(g4807,g4473);
  not NOT_2748(I9236,g6939);
  not NOT_2749(g3967,I5223);
  not NOT_2750(I6561,g4707);
  not NOT_2751(g6588,I8632);
  not NOT_2752(I4935,g3369);
  not NOT_2753(I2596,g985);
  not NOT_2754(g6161,g5926);
  not NOT_2755(g1274,g856);
  not NOT_2756(g6361,I8147);
  not NOT_2757(g1426,I2445);
  not NOT_2758(g2196,I3337);
  not NOT_2759(I7600,g5605);
  not NOT_2760(g2803,g2440);
  not NOT_2761(I6004,g4159);
  not NOT_2762(g3229,I4486);
  not NOT_2763(I6986,g5230);
  not NOT_2764(g6051,g5824);
  not NOT_2765(g5270,I6927);
  not NOT_2766(g804,I1871);
  not NOT_2767(I3255,g1650);
  not NOT_2768(g2538,I3656);
  not NOT_2769(g1325,I2330);
  not NOT_2770(g1821,I2883);
  not NOT_2771(g844,g578);
  not NOT_2772(I3481,g1461);
  not NOT_2773(I8034,g6242);
  not NOT_2774(g4142,I5508);
  not NOT_2775(g4248,I5696);
  not NOT_2776(g2509,I3635);
  not NOT_2777(I6546,g4692);
  not NOT_2778(I3726,g2030);
  not NOT_2779(g4815,I6495);
  not NOT_2780(I5644,g4059);
  not NOT_2781(I8147,g6182);
  not NOT_2782(g5124,I6780);
  not NOT_2783(g6103,I7805);
  not NOT_2784(I5119,g3714);
  not NOT_2785(g4692,I6280);
  not NOT_2786(g2467,I3599);
  not NOT_2787(I8681,g6566);
  not NOT_2788(g4726,I6352);
  not NOT_2789(g5469,I7153);
  not NOT_2790(g4154,I5548);
  not NOT_2791(I2601,g1161);
  not NOT_2792(g6696,I8806);
  not NOT_2793(g1636,I2593);
  not NOT_2794(g3921,g3512);
  not NOT_2795(g5540,I7284);
  not NOT_2796(I5577,g4022);
  not NOT_2797(g1106,I2128);
  not NOT_2798(g6732,I8888);
  not NOT_2799(g853,g642);
  not NOT_2800(g2256,I3395);
  not NOT_2801(g1790,I2842);
  not NOT_2802(I2922,g1774);
  not NOT_2803(g6508,I8444);
  not NOT_2804(I5893,g3747);
  not NOT_2805(I3979,g1836);
  not NOT_2806(I2581,g946);
  not NOT_2807(I3112,g1439);
  not NOT_2808(g1461,I2460);
  not NOT_2809(g3462,g2679);
  not NOT_2810(g1756,I2779);
  not NOT_2811(g2381,I3528);
  not NOT_2812(I6789,g4871);
  not NOT_2813(g4783,I6441);
  not NOT_2814(g6043,g5824);
  not NOT_2815(I7871,g6097);
  not NOT_2816(I2460,g952);
  not NOT_2817(I3001,g1267);
  not NOT_2818(g4112,I5418);
  not NOT_2819(g4218,I5640);
  not NOT_2820(g2197,I3340);
  not NOT_2821(g4267,I5720);
  not NOT_2822(I4166,g2390);
  not NOT_2823(g2397,I3540);
  not NOT_2824(I4366,g2244);
  not NOT_2825(g5199,I6867);
  not NOT_2826(g5399,I7065);
  not NOT_2827(g1046,g489);
  not NOT_2828(I3761,g2505);
  not NOT_2829(g3788,g3466);
  not NOT_2830(g6034,g5824);
  not NOT_2831(g6434,I8300);
  not NOT_2832(g6565,I8579);
  not NOT_2833(I6299,g4438);
  not NOT_2834(g4293,I5750);
  not NOT_2835(g4129,I5469);
  not NOT_2836(g5797,I7596);
  not NOT_2837(I3830,g2179);
  not NOT_2838(I2995,g1742);
  not NOT_2839(g6147,I7871);
  not NOT_2840(g1345,I2382);
  not NOT_2841(g1841,I2929);
  not NOT_2842(g6347,I8103);
  not NOT_2843(I1832,g143);
  not NOT_2844(I2479,g1049);
  not NOT_2845(I7339,g5540);
  not NOT_2846(g1191,g38);
  not NOT_2847(I2668,g1011);
  not NOT_2848(g1391,I2424);
  not NOT_2849(I1853,g211);
  not NOT_2850(g3192,I4429);
  not NOT_2851(g6533,I8515);
  not NOT_2852(g3085,I4324);
  not NOT_2853(I3746,g2035);
  not NOT_2854(I7838,g5947);
  not NOT_2855(g4727,I6355);
  not NOT_2856(I4964,g3673);
  not NOT_2857(g3485,g2986);
  not NOT_2858(I2190,g297);
  not NOT_2859(g1695,g1106);
  not NOT_2860(g6697,I8809);
  not NOT_2861(g1637,I2596);
  not NOT_2862(g1107,I2131);
  not NOT_2863(g2631,I3773);
  not NOT_2864(g6596,I8656);
  not NOT_2865(g3854,I5071);
  not NOT_2866(I5106,g3247);
  not NOT_2867(I8597,g6445);
  not NOT_2868(g2817,g2461);
  not NOT_2869(I6244,g4519);
  not NOT_2870(I7077,g5281);
  not NOT_2871(g4703,I6299);
  not NOT_2872(g6413,I8249);
  not NOT_2873(I5790,g3803);
  not NOT_2874(g1858,I2964);
  not NOT_2875(I6078,g4387);
  not NOT_2876(I6340,g4561);
  not NOT_2877(I7643,g5752);
  not NOT_2878(I3068,g1439);
  not NOT_2879(g5923,I7701);
  not NOT_2880(I9038,g6833);
  not NOT_2881(I3468,g1802);
  not NOT_2882(I4279,g2230);
  not NOT_2883(I5756,g3922);
  not NOT_2884(g6820,I8997);
  not NOT_2885(g4624,g4265);
  not NOT_2886(I6959,g5089);
  not NOT_2887(I5622,g3914);
  not NOT_2888(g3219,I4462);
  not NOT_2889(I5027,g3267);
  not NOT_2890(I4318,g2171);
  not NOT_2891(I7634,g5727);
  not NOT_2892(I5427,g3726);
  not NOT_2893(g3031,I4246);
  not NOT_2894(g1115,g40);
  not NOT_2895(g6117,g5880);
  not NOT_2896(g1315,I2296);
  not NOT_2897(g1811,I2864);
  not NOT_2898(g1642,g809);
  not NOT_2899(I8479,g6482);
  not NOT_2900(g2585,I3708);
  not NOT_2901(I7104,g5273);
  not NOT_2902(I5904,g3749);
  not NOT_2903(I8668,g6530);
  not NOT_2904(g5886,g5753);
  not NOT_2905(I8840,g6657);
  not NOT_2906(g2041,I3152);
  not NOT_2907(g6601,I8671);
  not NOT_2908(I5514,g3882);
  not NOT_2909(I3349,g1334);
  not NOT_2910(I2053,g684);
  not NOT_2911(g5114,I6756);
  not NOT_2912(I5403,g3970);
  not NOT_2913(g5314,I6972);
  not NOT_2914(I2453,g952);
  not NOT_2915(g1654,g878);
  not NOT_2916(g4716,I6330);
  not NOT_2917(g4149,I5529);
  not NOT_2918(g6922,I9203);
  not NOT_2919(I8156,g6167);
  not NOT_2920(I3198,g1819);
  not NOT_2921(I3855,g2550);
  not NOT_2922(I5391,g3975);
  not NOT_2923(g3911,I5148);
  not NOT_2924(g6581,g6493);
  not NOT_2925(g4848,I6552);
  not NOT_2926(I5637,g3914);
  not NOT_2927(g1880,g1603);
  not NOT_2928(g4198,I5618);
  not NOT_2929(g4699,I6289);
  not NOT_2930(g6597,I8659);
  not NOT_2931(g4855,I6573);
  not NOT_2932(g4398,I5893);
  not NOT_2933(g2772,I3961);
  not NOT_2934(I4321,g1917);
  not NOT_2935(g5136,I6786);
  not NOT_2936(g3225,I4474);
  not NOT_2937(I5223,g3537);
  not NOT_2938(g2743,g2333);
  not NOT_2939(g6784,I8940);
  not NOT_2940(g2890,g1875);
  not NOT_2941(g3073,I4300);
  not NOT_2942(g1978,g1387);
  not NOT_2943(g3796,g3388);
  not NOT_2944(g1017,I2053);
  not NOT_2945(I2929,g1659);
  not NOT_2946(g798,I1868);
  not NOT_2947(g2505,I3629);
  not NOT_2948(I3644,g1685);
  not NOT_2949(g3124,I4371);
  not NOT_2950(g1935,I3040);
  not NOT_2951(g3980,I5264);
  not NOT_2952(g2856,g2010);
  not NOT_2953(g2734,I3902);
  not NOT_2954(I8432,g6411);
  not NOT_2955(I3319,g1636);
  not NOT_2956(g1982,I3093);
  not NOT_2957(g754,I1850);
  not NOT_2958(g4524,I6084);
  not NOT_2959(g836,g349);
  not NOT_2960(I8453,g6414);
  not NOT_2961(g6840,I9041);
  not NOT_2962(I4519,g2788);
  not NOT_2963(g4644,I6231);
  not NOT_2964(I3152,g1322);
  not NOT_2965(I3258,g1760);
  not NOT_2966(g3540,I4762);
  not NOT_2967(I3352,g1285);
  not NOT_2968(g1328,I2337);
  not NOT_2969(g5887,g5742);
  not NOT_2970(g4119,I5439);
  not NOT_2971(g5465,I7143);
  not NOT_2972(g1542,g878);
  not NOT_2973(g1330,I2343);
  not NOT_2974(g3177,I4414);
  not NOT_2975(I3717,g2154);
  not NOT_2976(g5230,I6895);
  not NOT_2977(g845,g582);
  not NOT_2978(g4152,I5542);
  not NOT_2979(g6501,I8423);
  not NOT_2980(g4577,g4202);
  not NOT_2981(g4717,g4465);
  not NOT_2982(g5433,I7107);
  not NOT_2983(I5654,g3742);
  not NOT_2984(I6930,g5017);
  not NOT_2985(g2863,g2296);
  not NOT_2986(I6464,g4562);
  not NOT_2987(I3599,g1484);
  not NOT_2988(g2713,I3868);
  not NOT_2989(I3274,g1773);
  not NOT_2990(g4386,I5865);
  not NOT_2991(g3199,g1861);
  not NOT_2992(g5550,g5331);
  not NOT_2993(I3614,g1295);
  not NOT_2994(g3781,I4976);
  not NOT_2995(I3370,g1805);
  not NOT_2996(g5137,I6789);
  not NOT_2997(g5395,I7061);
  not NOT_2998(g5891,g5731);
  not NOT_2999(g3898,g3575);
  not NOT_3000(g3900,g3575);
  not NOT_3001(I3325,g1340);
  not NOT_3002(g4426,I5929);
  not NOT_3003(I2735,g1118);
  not NOT_3004(g3797,g3388);
  not NOT_3005(I9085,g6850);
  not NOT_3006(g1902,I3001);
  not NOT_3007(g6163,g5926);
  not NOT_3008(g4614,g4308);
  not NOT_3009(I2782,g1177);
  not NOT_3010(I7679,g5726);
  not NOT_3011(g6363,I8153);
  not NOT_3012(g4370,I5831);
  not NOT_3013(I8626,g6543);
  not NOT_3014(g3510,g2709);
  not NOT_3015(I5612,g3910);
  not NOT_3016(g6032,g5770);
  not NOT_3017(g4125,I5457);
  not NOT_3018(g2688,I3836);
  not NOT_3019(g2857,I4059);
  not NOT_3020(g3291,g3037);
  not NOT_3021(I3083,g1426);
  not NOT_3022(g2976,g2197);
  not NOT_3023(g1823,I2887);
  not NOT_3024(I2949,g1263);
  not NOT_3025(g1366,I2402);
  not NOT_3026(g5266,I6923);
  not NOT_3027(I2627,g1053);
  not NOT_3028(g1056,g89);
  not NOT_3029(g6568,I8588);
  not NOT_3030(I5328,g3502);
  not NOT_3031(g1529,g1076);
  not NOT_3032(I7805,g5923);
  not NOT_3033(I5542,g3984);
  not NOT_3034(I2998,g1257);
  not NOT_3035(g1649,g985);
  not NOT_3036(g1348,I2385);
  not NOT_3037(g3259,g2996);
  not NOT_3038(I4358,g2525);
  not NOT_3039(g5248,g4911);
  not NOT_3040(g4636,g4286);
  not NOT_3041(g1355,I2394);
  not NOT_3042(g4106,I5400);
  not NOT_3043(g5255,g4933);
  not NOT_3044(g3852,I5065);
  not NOT_3045(I9031,g6809);
  not NOT_3046(g2760,I3942);
  not NOT_3047(g3488,g2728);
  not NOT_3048(I8894,g6709);
  not NOT_3049(g4790,I6456);
  not NOT_3050(g5692,I7451);
  not NOT_3051(I4587,g2962);
  not NOT_3052(g5097,I6733);
  not NOT_3053(g5726,I7487);
  not NOT_3054(g4187,I5591);
  not NOT_3055(I9176,g6881);
  not NOT_3056(g4387,I5868);
  not NOT_3057(I9005,g6817);
  not NOT_3058(g1063,g675);
  not NOT_3059(g3886,g3346);
  not NOT_3060(g4622,g4252);
  not NOT_3061(g2608,I3746);
  not NOT_3062(I2919,g1787);
  not NOT_3063(g2779,g2394);
  not NOT_3064(g4904,g4812);
  not NOT_3065(g3114,I4362);
  not NOT_3066(I2952,g1594);
  not NOT_3067(g1279,g848);
  not NOT_3068(g4514,I6054);
  not NOT_3069(g1720,g1111);
  not NOT_3070(g4003,g3441);
  not NOT_3071(g1118,g36);
  not NOT_3072(I3391,g1646);
  not NOT_3073(g1318,I2309);
  not NOT_3074(g4403,I5904);
  not NOT_3075(I5490,g3832);
  not NOT_3076(g5112,I6750);
  not NOT_3077(g2588,I3717);
  not NOT_3078(g4145,I5517);
  not NOT_3079(g4841,I6531);
  not NOT_3080(I8603,g6449);
  not NOT_3081(g2361,I3513);
  not NOT_3082(I6769,g4786);
  not NOT_3083(g4763,I6397);
  not NOT_3084(g4191,I5603);
  not NOT_3085(g4391,I5876);
  not NOT_3086(I5056,g3567);
  not NOT_3087(I2986,g1504);
  not NOT_3088(I3307,g1339);
  not NOT_3089(g1193,I2204);
  not NOT_3090(I5529,g3854);
  not NOT_3091(I4420,g2096);
  not NOT_3092(I5148,g3450);
  not NOT_3093(g3136,I4382);
  not NOT_3094(g2327,I3481);
  not NOT_3095(I6918,g5124);
  not NOT_3096(I4507,g2739);
  not NOT_3097(g5329,I6989);
  not NOT_3098(g1549,g878);
  not NOT_3099(g4107,I5403);
  not NOT_3100(I7042,g5310);
  not NOT_3101(g947,g74);
  not NOT_3102(g6894,I9149);
  not NOT_3103(g1834,I2916);
  not NOT_3104(I4794,g2814);
  not NOT_3105(g4307,I5774);
  not NOT_3106(I5851,g3739);
  not NOT_3107(g4536,I6118);
  not NOT_3108(I3858,g2197);
  not NOT_3109(I8702,g6572);
  not NOT_3110(g2346,I3496);
  not NOT_3111(g6735,I8897);
  not NOT_3112(I3016,g1754);
  not NOT_3113(I2970,g1504);
  not NOT_3114(g5727,I7490);
  not NOT_3115(I7164,g5433);
  not NOT_3116(g2103,I3225);
  not NOT_3117(g858,g301);
  not NOT_3118(I2925,g1762);
  not NOT_3119(g4858,I6582);
  not NOT_3120(I3522,g1664);
  not NOT_3121(g4016,I5320);
  not NOT_3122(I3115,g1519);
  not NOT_3123(I3251,g1471);
  not NOT_3124(I3811,g2145);
  not NOT_3125(I8276,g6303);
  not NOT_3126(g1321,I2318);
  not NOT_3127(I3047,g1426);
  not NOT_3128(g1670,I2648);
  not NOT_3129(g3228,I4483);
  not NOT_3130(g3465,g2986);
  not NOT_3131(g3322,g3070);
  not NOT_3132(I5463,g3783);
  not NOT_3133(g3230,I4489);
  not NOT_3134(g4522,I6078);
  not NOT_3135(g4115,I5427);
  not NOT_3136(g2753,I3927);
  not NOT_3137(g4251,I5705);
  not NOT_3138(g1232,I2228);
  not NOT_3139(I4300,g2234);
  not NOT_3140(g6526,I8494);
  not NOT_3141(g1813,I2870);
  not NOT_3142(I8527,g6440);
  not NOT_3143(I8647,g6528);
  not NOT_3144(I2617,g1193);
  not NOT_3145(I5720,g4022);
  not NOT_3146(g2043,I3158);
  not NOT_3147(g6039,g5824);
  not NOT_3148(I8764,g6564);
  not NOT_3149(g2443,I3578);
  not NOT_3150(g6484,g6361);
  not NOT_3151(g3096,I4343);
  not NOT_3152(g5468,I7150);
  not NOT_3153(g1519,I2491);
  not NOT_3154(g1740,g1116);
  not NOT_3155(I7012,g5316);
  not NOT_3156(g6850,I9077);
  not NOT_3157(I6895,g5010);
  not NOT_3158(I1835,g205);
  not NOT_3159(g3845,I5050);
  not NOT_3160(I5843,g3851);
  not NOT_3161(g2316,I3468);
  not NOT_3162(I3537,g1305);
  not NOT_3163(I8503,g6434);
  not NOT_3164(g1552,g1030);
  not NOT_3165(I5457,g3766);
  not NOT_3166(g2565,I3675);
  not NOT_3167(g6583,I8617);
  not NOT_3168(g850,g602);
  not NOT_3169(g5576,g5415);
  not NOT_3170(g4537,g4410);
  not NOT_3171(I7029,g5149);
  not NOT_3172(g2347,I3499);
  not NOT_3173(I5686,g3942);
  not NOT_3174(I4123,g2043);
  not NOT_3175(g3807,I5006);
  not NOT_3176(g1586,g1052);
  not NOT_3177(g3859,I5078);
  not NOT_3178(g6276,I7960);
  not NOT_3179(g4612,g4320);
  not NOT_3180(g2914,g1928);
  not NOT_3181(g6616,I8710);
  not NOT_3182(I3629,g1759);
  not NOT_3183(g6561,I8567);
  not NOT_3184(I3328,g1273);
  not NOT_3185(I2738,g1236);
  not NOT_3186(I8617,g6539);
  not NOT_3187(g1341,I2376);
  not NOT_3188(g2413,I3553);
  not NOT_3189(I4351,g2233);
  not NOT_3190(g3342,g3086);
  not NOT_3191(g4128,I5466);
  not NOT_3192(g1710,g1109);
  not NOT_3193(g4629,g4276);
  not NOT_3194(I6485,g4603);
  not NOT_3195(g6527,I8497);
  not NOT_3196(g6404,I8226);
  not NOT_3197(g4328,g4092);
  not NOT_3198(I2140,g28);
  not NOT_3199(g1645,I2614);
  not NOT_3200(I2340,g1142);
  not NOT_3201(g4130,I5472);
  not NOT_3202(I5938,g4351);
  not NOT_3203(I7963,g6276);
  not NOT_3204(I3800,g2145);
  not NOT_3205(g3481,g2612);
  not NOT_3206(I2907,g1498);
  not NOT_3207(g2820,g2470);
  not NOT_3208(g2936,g2026);
  not NOT_3209(g5524,I7264);
  not NOT_3210(g6503,I8429);
  not NOT_3211(g3354,g3096);
  not NOT_3212(I4410,g2088);
  not NOT_3213(I7808,g5919);
  not NOT_3214(g2117,I3244);
  not NOT_3215(g3960,I5204);
  not NOT_3216(g2317,I3471);
  not NOT_3217(g5119,I6769);
  not NOT_3218(g6925,I9208);
  not NOT_3219(I7707,g5701);
  not NOT_3220(I5606,g3821);
  not NOT_3221(g1659,I2638);
  not NOT_3222(g1358,g1119);
  not NOT_3223(g5352,I7002);
  not NOT_3224(g5577,g5420);
  not NOT_3225(g4213,I5633);
  not NOT_3226(g5717,I7478);
  not NOT_3227(I3902,g2576);
  not NOT_3228(g6120,I7832);
  not NOT_3229(g2922,g1960);
  not NOT_3230(g1587,g1123);
  not NOT_3231(I6812,g5110);
  not NOT_3232(I8991,g6788);
  not NOT_3233(g3783,I4980);
  not NOT_3234(g1111,I2143);
  not NOT_3235(I3090,g1504);
  not NOT_3236(I9008,g6818);
  not NOT_3237(g5893,g5753);
  not NOT_3238(g1275,g842);
  not NOT_3239(g6277,I7963);
  not NOT_3240(g2581,I3694);
  not NOT_3241(I3823,g2125);
  not NOT_3242(g3267,g3030);
  not NOT_3243(I4667,g2908);
  not NOT_3244(g3312,I4587);
  not NOT_3245(I7865,g6095);
  not NOT_3246(I4343,g2525);
  not NOT_3247(g2060,g1369);
  not NOT_3248(g6617,I8713);
  not NOT_3249(g6906,I9185);
  not NOT_3250(g5975,g5821);
  not NOT_3251(g4512,I6048);
  not NOT_3252(I4282,g2525);
  not NOT_3253(g2460,I3590);
  not NOT_3254(I7604,g5605);
  not NOT_3255(I8907,g6702);
  not NOT_3256(I3056,g1519);
  not NOT_3257(g3001,I4198);
  not NOT_3258(g1174,g37);
  not NOT_3259(g4823,I6507);
  not NOT_3260(I2663,g1006);
  not NOT_3261(g4166,I5568);
  not NOT_3262(g6516,g6409);
  not NOT_3263(g5274,I6933);
  not NOT_3264(I8435,g6413);
  not NOT_3265(I3148,g1595);
  not NOT_3266(I8690,g6571);
  not NOT_3267(g1985,I3096);
  not NOT_3268(I4334,g2256);
  not NOT_3269(I8482,g6461);
  not NOT_3270(g2739,I3906);
  not NOT_3271(g3761,g3605);
  not NOT_3272(I3155,g1612);
  not NOT_3273(I3355,g1608);
  not NOT_3274(I2402,g774);
  not NOT_3275(g4529,I6099);
  not NOT_3276(g1284,g851);
  not NOT_3277(g4148,I5526);
  not NOT_3278(I6733,g4773);
  not NOT_3279(I8656,g6532);
  not NOT_3280(g3830,I5019);
  not NOT_3281(I9122,g6864);
  not NOT_3282(g2079,g1348);
  not NOT_3283(g4155,I5551);
  not NOT_3284(g4851,I6561);
  not NOT_3285(g6892,I9143);
  not NOT_3286(g1832,I2910);
  not NOT_3287(I9230,g6936);
  not NOT_3288(g1853,I2955);
  not NOT_3289(g2840,g2538);
  not NOT_3290(I2877,g1123);
  not NOT_3291(I5879,g3745);
  not NOT_3292(g5544,g5331);
  not NOT_3293(g2390,I3531);
  not NOT_3294(I6324,g4450);
  not NOT_3295(g1559,g965);
  not NOT_3296(I6069,g4213);
  not NOT_3297(I8110,g6143);
  not NOT_3298(g4463,g4364);
  not NOT_3299(g943,g496);
  not NOT_3300(g1931,I3034);
  not NOT_3301(g6709,I8837);
  not NOT_3302(g3932,I5169);
  not NOT_3303(I6540,g4714);
  not NOT_3304(I3720,g2155);
  not NOT_3305(g6078,g5801);
  not NOT_3306(I1871,g281);
  not NOT_3307(I6377,g4569);
  not NOT_3308(g5061,I6701);
  not NOT_3309(g6478,I8342);
  not NOT_3310(I2464,g850);
  not NOT_3311(I3367,g1283);
  not NOT_3312(g5387,I7051);
  not NOT_3313(I9137,g6864);
  not NOT_3314(g1905,I3004);
  not NOT_3315(I8002,g6110);
  not NOT_3316(g866,g314);
  not NOT_3317(I2785,g1222);
  not NOT_3318(I7086,g5281);
  not NOT_3319(I5615,g3914);
  not NOT_3320(g6035,g5824);
  not NOT_3321(g4720,I6340);
  not NOT_3322(I3843,g2145);
  not NOT_3323(g4118,I5436);
  not NOT_3324(g4619,g4248);
  not NOT_3325(g6517,I8467);
  not NOT_3326(g1204,g39);
  not NOT_3327(g3677,g3140);
  not NOT_3328(g6876,I9095);
  not NOT_3329(g4843,I6537);
  not NOT_3330(g3866,I5091);
  not NOT_3331(g2954,g2381);
  not NOT_3332(I4593,g2966);
  not NOT_3333(g5046,I6680);
  not NOT_3334(g2163,I3288);
  not NOT_3335(g6656,I8764);
  not NOT_3336(g4193,I5609);
  not NOT_3337(I2237,g465);
  not NOT_3338(g2032,g1749);
  not NOT_3339(g4393,I5882);
  not NOT_3340(I5545,g3814);
  not NOT_3341(g5403,I7069);
  not NOT_3342(I1838,g206);
  not NOT_3343(g3848,I5059);
  not NOT_3344(I5591,g3821);
  not NOT_3345(I4264,g2212);
  not NOT_3346(I2394,g719);
  not NOT_3347(g5391,I7055);
  not NOT_3348(g2568,I3678);
  not NOT_3349(I2731,g1117);
  not NOT_3350(I4050,g2059);
  not NOT_3351(g3241,I4522);
  not NOT_3352(g2912,g2001);
  not NOT_3353(g4121,I5445);
  not NOT_3354(g1969,I3080);
  not NOT_3355(I3232,g1782);
  not NOT_3356(g4321,I5790);
  not NOT_3357(g5307,I6959);
  not NOT_3358(g2157,I3278);
  not NOT_3359(g5536,g5467);
  not NOT_3360(g2357,I3509);
  not NOT_3361(g1123,I2165);
  not NOT_3362(g1323,I2324);
  not NOT_3363(g4625,g4267);
  not NOT_3364(I3909,g2044);
  not NOT_3365(g4232,I5674);
  not NOT_3366(g6402,I8220);
  not NOT_3367(g6824,I9005);
  not NOT_3368(g1666,g1088);
  not NOT_3369(g4938,I6630);
  not NOT_3370(I6819,g5019);
  not NOT_3371(g6236,g6070);
  not NOT_3372(I3519,g1305);
  not NOT_3373(I8295,g6295);
  not NOT_3374(I2955,g1729);
  not NOT_3375(I7487,g5684);
  not NOT_3376(g856,g654);
  not NOT_3377(I6923,g5124);
  not NOT_3378(g1528,g878);
  not NOT_3379(I5204,g3534);
  not NOT_3380(I5630,g3914);
  not NOT_3381(I6488,g4603);
  not NOT_3382(g1351,I2388);
  not NOT_3383(g1648,I2623);
  not NOT_3384(I2814,g1222);
  not NOT_3385(g1875,I2970);
  not NOT_3386(g4519,I6069);
  not NOT_3387(g5115,I6759);
  not NOT_3388(g6590,I8638);
  not NOT_3389(g5251,g5069);
  not NOT_3390(g6877,I9098);
  not NOT_3391(g3258,I4537);
  not NOT_3392(I4777,g2962);
  not NOT_3393(I6701,g4726);
  not NOT_3394(g5315,g5116);
  not NOT_3395(g3867,I5094);
  not NOT_3396(I2150,g10);
  not NOT_3397(g1655,g985);
  not NOT_3398(g6657,I8767);
  not NOT_3399(g4606,g4193);
  not NOT_3400(I3687,g1814);
  not NOT_3401(I8089,g6120);
  not NOT_3402(I2773,g1191);
  not NOT_3403(g5874,I7634);
  not NOT_3404(g1410,g1233);
  not NOT_3405(I8966,g6796);
  not NOT_3406(I5750,g4022);
  not NOT_3407(I7045,g5167);
  not NOT_3408(I6114,g4405);
  not NOT_3409(g3975,I5249);
  not NOT_3410(I7173,g5436);
  not NOT_3411(g1884,I2979);
  not NOT_3412(I7091,g5281);
  not NOT_3413(g6899,I9164);
  not NOT_3414(I4799,g2967);
  not NOT_3415(I2212,g123);
  not NOT_3416(g929,g49);
  not NOT_3417(g6785,I8943);
  not NOT_3418(g5880,g5824);
  not NOT_3419(I5040,g3271);
  not NOT_3420(I2967,g1682);
  not NOT_3421(g5537,g5385);
  not NOT_3422(g2778,g2391);
  not NOT_3423(I1862,g278);
  not NOT_3424(I3525,g1461);
  not NOT_3425(g3370,g3124);
  not NOT_3426(g2894,g1891);
  not NOT_3427(I7007,g5314);
  not NOT_3428(g1372,I2408);
  not NOT_3429(g4141,I5505);
  not NOT_3430(g6563,I8573);
  not NOT_3431(I6008,g4163);
  not NOT_3432(I3691,g1732);
  not NOT_3433(g4525,I6087);
  not NOT_3434(g1143,I2172);
  not NOT_3435(g3984,g3564);
  not NOT_3436(I8150,g6185);
  not NOT_3437(g1282,g849);
  not NOT_3438(I8438,g6416);
  not NOT_3439(g3083,I4318);
  not NOT_3440(g1988,I3099);
  not NOT_3441(I4802,g2877);
  not NOT_3442(I6972,g5135);
  not NOT_3443(g3483,g2716);
  not NOT_3444(I7261,g5458);
  not NOT_3445(g6194,I7906);
  not NOT_3446(g1334,I2355);
  not NOT_3447(I3158,g1829);
  not NOT_3448(I3659,g1491);
  not NOT_3449(I3358,g1323);
  not NOT_3450(g5328,I6986);
  not NOT_3451(I1927,g665);
  not NOT_3452(g6489,g6369);
  not NOT_3453(g5542,g5331);
  not NOT_3454(g5330,I6992);
  not NOT_3455(g3306,g3057);
  not NOT_3456(g2998,I4195);
  not NOT_3457(g4158,I5556);
  not NOT_3458(g4659,I6250);
  not NOT_3459(g1555,I2521);
  not NOT_3460(g3790,g3388);
  not NOT_3461(I3587,g1461);
  not NOT_3462(g1792,I2848);
  not NOT_3463(g2603,I3733);
  not NOT_3464(g2039,I3148);
  not NOT_3465(g3187,I4424);
  not NOT_3466(g2484,I3611);
  not NOT_3467(g3387,I4664);
  not NOT_3468(g3461,g2986);
  not NOT_3469(g4587,g4215);
  not NOT_3470(I6033,g4179);
  not NOT_3471(g5554,g5455);
  not NOT_3472(g3622,I4821);
  not NOT_3473(g4111,I5415);
  not NOT_3474(I8229,g6330);
  not NOT_3475(I9149,g6884);
  not NOT_3476(I2620,g1177);
  not NOT_3477(g1113,I2147);
  not NOT_3478(I4492,g3001);
  not NOT_3479(g4615,g4322);
  not NOT_3480(g2583,g1830);
  not NOT_3481(g3904,g3575);
  not NOT_3482(g3200,I4437);
  not NOT_3483(I6096,g4397);
  not NOT_3484(g3046,I4267);
  not NOT_3485(g899,I1924);
  not NOT_3486(g4374,I5837);
  not NOT_3487(I3284,g1702);
  not NOT_3488(g2919,g1937);
  not NOT_3489(g1908,I3007);
  not NOT_3490(I2788,g1236);
  not NOT_3491(g1094,I2122);
  not NOT_3492(I5618,g3821);
  not NOT_3493(g2952,g2381);
  not NOT_3494(I6337,g4455);
  not NOT_3495(I5343,g3599);
  not NOT_3496(g2276,I3425);
  not NOT_3497(g1567,I2537);
  not NOT_3498(g4284,I5739);
  not NOT_3499(g5512,I7254);
  not NOT_3500(g4545,g4416);
  not NOT_3501(g5090,g4741);
  not NOT_3502(g6409,g6285);
  not NOT_3503(g5490,I7190);
  not NOT_3504(I7689,g5708);
  not NOT_3505(g4380,I5851);
  not NOT_3506(I2842,g1177);
  not NOT_3507(g1776,I2821);
  not NOT_3508(g1593,g1054);
  not NOT_3509(g2004,I3115);
  not NOT_3510(g4853,I6567);
  not NOT_3511(g6836,I9031);
  not NOT_3512(I2485,g766);
  not NOT_3513(I3794,g2044);
  not NOT_3514(g2986,g2010);
  not NOT_3515(g4020,I5324);
  not NOT_3516(g6212,I7910);
  not NOT_3517(I5548,g4059);
  not NOT_3518(g5456,g5300);
  not NOT_3519(g2647,I3791);
  not NOT_3520(I8837,g6665);
  not NOT_3521(g5148,I6812);
  not NOT_3522(g5649,I7404);
  not NOT_3523(g4507,I6033);
  not NOT_3524(g3223,I4468);
  not NOT_3525(I4623,g2962);
  not NOT_3526(I1947,g699);
  not NOT_3527(g2764,g2357);
  not NOT_3528(I8620,g6541);
  not NOT_3529(I8462,g6430);
  not NOT_3530(I9119,g6855);
  not NOT_3531(I2854,g1236);
  not NOT_3532(g4559,g4187);
  not NOT_3533(g5155,g5099);
  not NOT_3534(g5355,I7007);
  not NOT_3535(I9152,g6889);
  not NOT_3536(g3016,I4223);
  not NOT_3537(g6229,g6036);
  not NOT_3538(g1160,I2179);
  not NOT_3539(g5260,g4938);
  not NOT_3540(I6081,g4388);
  not NOT_3541(I4375,g2254);
  not NOT_3542(g6822,g6786);
  not NOT_3543(g1641,I2604);
  not NOT_3544(g3251,I4534);
  not NOT_3545(I6692,g4720);
  not NOT_3546(g1450,I2453);
  not NOT_3547(g5063,g4799);
  not NOT_3548(I7910,g5905);
  not NOT_3549(I8249,g6289);
  not NOT_3550(g4628,g4273);
  not NOT_3551(g4515,I6057);
  not NOT_3552(g2120,I3251);
  not NOT_3553(I4285,g2555);
  not NOT_3554(g2320,I3474);
  not NOT_3555(g4100,I5382);
  not NOT_3556(g1724,I2724);
  not NOT_3557(g3874,I5103);
  not NOT_3558(I2958,g1257);
  not NOT_3559(I5094,g3705);
  not NOT_3560(I2376,g729);
  not NOT_3561(I8485,g6479);
  not NOT_3562(g5720,I7481);
  not NOT_3563(I2405,g1112);
  not NOT_3564(g2906,g1911);
  not NOT_3565(g2789,g2410);
  not NOT_3566(g1878,I2973);
  not NOT_3567(g5118,I6766);
  not NOT_3568(I9170,g6883);
  not NOT_3569(I1917,g48);
  and AND2_0(g2771,g2497,g1975);
  and AND2_1(g6620,g6516,g6117);
  and AND2_2(g5193,g532,g4967);
  and AND4_0(I5360,g3532,g3536,g3539,g3544);
  and AND2_3(g5598,g5046,g5509);
  and AND2_4(g6249,g1332,g5892);
  and AND2_5(g4666,g4630,g4627);
  and AND2_6(g3629,g2809,g2738);
  and AND2_7(g3328,g2701,g1894);
  and AND2_8(g6085,g1161,g5731);
  and AND2_9(g4351,g166,g3776);
  and AND2_10(g4648,g4407,g79);
  and AND2_11(g5232,g548,g4980);
  and AND2_12(g2340,g1398,g1387);
  and AND2_13(g5938,g5114,g5791);
  and AND2_14(g5909,g5787,g3384);
  and AND2_15(g1802,g89,g1064);
  and AND2_16(g3554,g2941,g179);
  and AND2_17(g4410,g3903,g1474);
  and AND2_18(g6640,g1612,g6549);
  and AND2_19(g4172,g3930,g1366);
  and AND2_20(g4372,g406,g3790);
  and AND2_21(g3512,g2928,g1764);
  and AND2_22(g3490,g353,g2959);
  and AND2_23(g4667,g4653,g4651);
  and AND2_24(g3166,g2042,g1233);
  and AND2_25(g3366,g248,g2893);
  and AND2_26(g6829,g6806,g5958);
  and AND2_27(g3649,g3104,g2764);
  and AND2_28(g6911,g6904,g6902);
  and AND2_29(g3155,g248,g2461);
  and AND2_30(g3698,g2284,g2835);
  and AND2_31(g6270,g1726,g6062);
  and AND2_32(g4792,g1417,g4471);
  and AND3_0(g6473,g2036,g6397,g1628);
  and AND2_33(g4621,g3953,g4364);
  and AND2_34(g5158,g504,g4993);
  and AND2_35(g6124,g5705,g5958);
  and AND2_36(g6324,g3880,g6212);
  and AND3_1(g6469,g2121,g2032,g6394);
  and AND2_37(g3279,g2599,g2612);
  and AND2_38(g3619,g2449,g3057);
  and AND2_39(g3167,g1883,g921);
  and AND2_40(g5311,g5013,g4468);
  and AND2_41(g3367,g2809,g1960);
  and AND2_42(g3652,g2544,g3096);
  and AND3_2(g3843,g2856,g945,g3533);
  and AND2_43(g4593,g4277,g947);
  and AND2_44(g3686,g2256,g2819);
  and AND2_45(g5180,g414,g4950);
  and AND2_46(g5380,g188,g5264);
  and AND2_47(g4160,g3923,g1345);
  and AND2_48(g3321,g2252,g2713);
  and AND2_49(g2089,g1123,g1578);
  and AND2_50(g6245,g1329,g5889);
  and AND2_51(g4360,g184,g3785);
  and AND2_52(g3670,g2234,g2792);
  and AND2_53(g3625,g2619,g2320);
  and AND2_54(g6291,g5210,g6161);
  and AND2_55(g4050,I5359,I5360);
  and AND2_56(g5559,g5024,g5453);
  and AND2_57(g6144,g3183,g5997);
  and AND2_58(g6344,g6272,g6080);
  and AND2_59(g2948,g2137,g1595);
  and AND2_60(g6259,g1699,g6044);
  and AND2_61(g4179,g390,g3902);
  and AND2_62(g2955,g2381,g297);
  and AND2_63(g6088,g1143,g5753);
  and AND2_64(g6852,g6847,g2295);
  and AND2_65(g6923,g6918,g6917);
  and AND2_66(g5515,g590,g5364);
  and AND2_67(g1499,g1101,g1094);
  and AND2_68(g4835,g4533,g4530);
  and AND2_69(g3687,g2245,g2820);
  and AND3_3(g4271,g2121,g1749,g4004);
  and AND3_4(g4611,g3985,g119,g4300);
  and AND2_70(g3341,g2998,g2709);
  and AND2_71(g6650,g6580,g6235);
  and AND2_72(g4541,g631,g4199);
  and AND2_73(g3645,g2497,g3090);
  and AND2_74(g5123,g4670,g1936);
  and AND2_75(g3691,g2268,g2828);
  and AND2_76(g4209,g3816,g865);
  and AND2_77(g4353,g3989,g3332);
  and AND2_78(g6336,g6246,g6065);
  and AND2_79(g6768,g6750,g3477);
  and AND2_80(g4744,g3434,g4582);
  and AND2_81(g3659,g2672,g2361);
  and AND2_82(g5351,g5326,g3459);
  and AND2_83(g3358,g2842,g1369);
  and AND2_84(g5648,g4507,g5545);
  and AND2_85(g6934,g6932,g3605);
  and AND2_86(g3275,g2172,g2615);
  and AND2_87(g3311,g218,g2872);
  and AND2_88(g5410,g378,g5274);
  and AND2_89(g3615,g2422,g3046);
  and AND2_90(g2062,g1499,g1666);
  and AND2_91(g3374,g2809,g1969);
  and AND2_92(g4600,g4054,g4289);
  and AND2_93(g6096,g1193,g5753);
  and AND2_94(g1436,g834,g830);
  and AND2_95(g5172,g441,g4877);
  and AND2_96(g3180,g260,g2506);
  and AND2_97(g5618,g5506,g4933);
  and AND2_98(g5143,g157,g5099);
  and AND2_99(g6913,g6900,g6898);
  and AND2_100(g5235,g554,g4980);
  and AND2_101(g4580,g706,g4262);
  and AND2_102(g2085,g1123,g1567);
  and AND2_103(g6266,g1721,g6057);
  and AND2_104(g5555,g5014,g5442);
  and AND2_105(g2941,g2166,g170);
  and AND2_106(g6248,g465,g5894);
  and AND2_107(g6342,g6264,g6076);
  and AND2_108(g5621,g5508,g4943);
  and AND2_109(g3628,g2449,g3070);
  and AND2_110(g6255,g1335,g5895);
  and AND2_111(g6081,g1177,g5731);
  and AND2_112(g3630,g3167,g1756);
  and AND2_113(g6692,g6616,g6615);
  and AND2_114(g3300,g2232,g2682);
  and AND2_115(g6154,g3219,g6015);
  and AND2_116(g6354,g5866,g6193);
  and AND2_117(g4184,g3934,g2136);
  and AND2_118(g5494,g5443,g3455);
  and AND2_119(g4384,g414,g3797);
  and AND2_120(g4339,g3971,g3289);
  and AND2_121(g4838,g4648,g84);
  and AND2_122(g3123,g230,g2391);
  and AND2_123(g3323,g2253,g2716);
  and AND2_124(g4672,g4635,g4631);
  and AND2_125(g2733,g2422,g1943);
  and AND2_126(g3666,g3128,g2787);
  and AND2_127(g6129,g5717,g5975);
  and AND2_128(g6329,g3888,g6212);
  and AND2_129(g2073,g1088,g1499);
  and AND2_130(g5360,g4431,g5160);
  and AND2_131(g6828,g6803,g5958);
  and AND2_132(g5050,g4285,g4807);
  and AND2_133(g3351,g2760,g1931);
  and AND2_134(g6830,g6809,g5975);
  and AND2_135(g3648,g2722,g2343);
  and AND2_136(g3655,g2197,g2768);
  and AND3_5(g1706,g766,g719,g729);
  and AND2_137(g6068,g5824,g1726);
  and AND2_138(g4044,g410,g3388);
  and AND3_6(g6468,g2032,g6394,g1609);
  and AND2_139(g3172,g2449,g2491);
  and AND2_140(g3278,g2175,g2628);
  and AND2_141(g3372,g254,g2905);
  and AND2_142(g2781,g2544,g1982);
  and AND2_143(g3618,g3016,g2712);
  and AND2_144(g3667,g2245,g2789);
  and AND2_145(g3143,g242,g2437);
  and AND2_146(g3282,g131,g2863);
  and AND2_147(g6716,g6682,g932);
  and AND2_148(g6149,g3200,g5997);
  and AND2_149(g3693,g2256,g2830);
  and AND2_150(g3134,g230,g2413);
  and AND2_151(g3334,g236,g2883);
  and AND3_7(g6848,g3741,g328,g6843);
  and AND2_152(g5153,g492,g4904);
  and AND2_153(g5209,g560,g5025);
  and AND2_154(g5353,g5327,g3463);
  and AND2_155(g6241,g1325,g5887);
  and AND2_156(g1808,g706,g49);
  and AND2_157(g3113,g224,g2364);
  and AND2_158(g5558,g5018,g5450);
  and AND2_159(g6644,g6575,g6230);
  and AND2_160(g6152,g3212,g6015);
  and AND2_161(g6258,g512,g5899);
  and AND2_162(g4178,g3959,g2110);
  and AND2_163(g1575,g980,g965);
  and AND2_164(g4378,g410,g3792);
  and AND2_165(g4831,g4528,g4524);
  and AND2_166(g4182,g394,g3904);
  and AND2_167(g5492,g5441,g3452);
  and AND2_168(g5600,g5502,g4900);
  and AND2_169(g6614,g932,g6556);
  and AND2_170(g4947,g184,g4741);
  and AND2_171(g3360,g2783,g1947);
  and AND2_172(g6125,g5708,g5975);
  and AND2_173(g1419,g613,g918);
  and AND2_174(g3641,g2644,g2333);
  and AND2_175(g4873,g4838,g4173);
  and AND2_176(g4037,g2896,g3388);
  and AND2_177(g3724,g117,g3251);
  and AND2_178(g4495,g3913,g4292);
  and AND2_179(g3379,g3104,g1988);
  and AND2_180(g5175,g5094,g1384);
  and AND2_181(g3658,g3118,g2776);
  and AND2_182(g6061,g5824,g1711);
  and AND2_183(g5500,g5430,g5074);
  and AND2_184(g3611,g2370,g3037);
  and AND2_185(g2137,g760,g1638);
  and AND2_186(g4042,g406,g3388);
  and AND2_187(g5184,g453,g4877);
  and AND2_188(g4442,g4239,g2882);
  and AND2_189(g4164,g3958,g2091);
  and AND2_190(g2807,g2568,g2001);
  and AND2_191(g5424,g390,g5296);
  and AND2_192(g6145,g3187,g6015);
  and AND2_193(g2859,g2112,g1649);
  and AND3_8(g3997,g1250,g3425,g2849);
  and AND2_194(g4054,g3694,g69);
  and AND2_195(g6345,g6273,g6083);
  and AND2_196(g3132,g2306,g1206);
  and AND2_197(g3680,g2245,g2805);
  and AND2_198(g6637,g1842,g6549);
  and AND2_199(g3353,g3162,g2921);
  and AND2_200(g2142,g1793,g1777);
  and AND2_201(g2255,g1706,g736);
  and AND2_202(g6159,g3177,g6015);
  and AND2_203(g2081,g1094,g1546);
  and AND2_204(g3558,g338,g3199);
  and AND2_205(g5499,g5451,g3462);
  and AND2_206(g4389,g449,g3798);
  and AND2_207(g4171,g3956,g2104);
  and AND2_208(g6315,g3849,g6194);
  and AND2_209(g4371,g461,g3789);
  and AND3_9(g4429,g923,g4253,g2936);
  and AND2_210(g4787,g2937,g4628);
  and AND2_211(g6047,g5824,g1692);
  and AND2_212(g6874,g6873,g2060);
  and AND2_213(g2267,g1716,g791);
  and AND3_10(g5444,g4545,g5256,g1574);
  and AND2_214(g5269,g557,g5025);
  and AND2_215(g1407,g301,g866);
  and AND2_216(g4684,g4584,g1341);
  and AND2_217(g4791,g3936,g4636);
  and AND2_218(g6243,g500,g5890);
  and AND2_219(g6935,g6933,g3622);
  and AND2_220(g2746,g2473,g1954);
  and AND2_221(g4759,g536,g4500);
  and AND2_222(g6128,g5590,g5958);
  and AND2_223(g5414,g382,g5278);
  and AND2_224(g6130,g5720,g5958);
  and AND2_225(g5660,g4509,g5549);
  and AND2_226(g3375,g260,g2912);
  and AND2_227(g4449,g4266,g2887);
  and AND2_228(g3651,g3064,g2766);
  and AND2_229(g4865,g4776,g1849);
  and AND2_230(g2953,g2381,g293);
  and AND2_231(g2068,g1541,g1546);
  and AND2_232(g3285,g2195,g2653);
  and AND2_233(g4833,g4521,g4516);
  and AND2_234(g5178,g516,g4993);
  and AND2_235(g5679,g74,g5576);
  and AND2_236(g5378,g179,g5260);
  and AND2_237(g3339,g2734,g1914);
  and AND2_238(g1689,g766,g719);
  and AND2_239(g5182,g520,g4993);
  and AND2_240(g2699,g2397,g1905);
  and AND2_241(g2747,g2449,g1957);
  and AND2_242(g6090,g1161,g5742);
  and AND2_243(g4362,g3996,g3355);
  and AND2_244(g3672,g3136,g2800);
  and AND2_245(g4052,g418,g3388);
  and AND2_246(g3643,g2518,g3086);
  and AND2_247(g4452,g3820,g4227);
  and AND2_248(g6056,g5824,g1699);
  and AND2_249(g1826,g714,g710);
  and AND2_250(g6148,g3196,g6015);
  and AND2_251(g6348,g5869,g6211);
  and AND2_252(g5560,g5044,g5456);
  and AND2_253(g3634,g2179,g2744);
  and AND2_254(g6155,g2588,g5997);
  and AND2_255(g6851,g6846,g2293);
  and AND2_256(g3551,g2937,g938);
  and AND2_257(g3099,g218,g2350);
  and AND2_258(g3304,g2857,g1513);
  and AND2_259(g4486,g716,g4195);
  and AND2_260(g3499,g357,g2961);
  and AND2_261(g4730,g1423,g4565);
  and AND2_262(g5632,g4494,g5538);
  and AND2_263(g5095,g4794,g951);
  and AND2_264(g6260,g1703,g6048);
  and AND2_265(g4185,g398,g3906);
  and AND2_266(g1609,g760,g754);
  and AND2_267(g5495,g5444,g3456);
  and AND4_1(g2577,g1743,g1797,g1793,g1138);
  and AND2_268(g3613,g2604,g2312);
  and AND2_269(g6619,g6515,g6115);
  and AND2_270(g6318,g3865,g6212);
  and AND4_2(g2026,g1359,g1402,g1398,g901);
  and AND2_271(g5164,g437,g4877);
  and AND2_272(g5364,g574,g5194);
  and AND2_273(g5233,g551,g4980);
  and AND2_274(g2821,g1890,g910);
  and AND2_275(g3729,g327,g3441);
  and AND2_276(g5454,g5256,g4549);
  and AND2_277(g5553,g5012,g5440);
  and AND2_278(g6321,g3873,g6212);
  and AND2_279(g3660,g2568,g3110);
  and AND3_11(g6625,g2121,g1595,g6538);
  and AND2_280(g4045,g3425,g123);
  and AND2_281(g4445,g4235,g1854);
  and AND2_282(g6253,g508,g5896);
  and AND2_283(g4373,g4001,g3370);
  and AND2_284(g5189,g528,g4993);
  and AND2_285(g4491,g3554,g4215);
  and AND2_286(g6909,g6896,g6894);
  and AND2_287(g4169,g3966,g2099);
  and AND2_288(g5171,g406,g4950);
  and AND2_289(g4369,g3999,g3364);
  and AND2_290(g3679,g2245,g2803);
  and AND2_291(g4602,g4407,g4293);
  and AND2_292(g5371,g152,g5248);
  and AND2_293(g3378,g3136,g2932);
  and AND2_294(g5429,g398,g5304);
  and AND2_295(g4407,g4054,g74);
  and AND2_296(g5956,g5783,g5425);
  and AND2_297(g4868,g4774,g2891);
  and AND2_298(g5675,g64,g5574);
  and AND2_299(g3135,g2370,g2416);
  and AND2_300(g4459,g4245,g1899);
  and AND2_301(g3335,g230,g2884);
  and AND2_302(g3831,g2330,g3425);
  and AND2_303(g3182,g2473,g2512);
  and AND2_304(g3288,g2631,g2634);
  and AND2_305(g3382,g3136,g2934);
  and AND2_306(g4793,g4277,g4639);
  and AND2_307(g4015,g445,g3388);
  and AND2_308(g2107,g1583,g1543);
  and AND2_309(g6141,g3173,g5997);
  and AND2_310(g6341,g6261,g6074);
  and AND2_311(g6645,g6576,g6231);
  and AND2_312(g3632,g3043,g2743);
  and AND2_313(g3437,g837,g2853);
  and AND2_314(g3653,g2215,g2767);
  and AND2_315(g5201,g4859,g5084);
  and AND2_316(g3208,g895,g2551);
  and AND2_317(g3302,g212,g2867);
  and AND2_318(g6158,g2594,g6015);
  and AND2_319(g5449,g4545,g5246);
  and AND2_320(g5604,g5059,g5521);
  and AND2_321(g5098,g4021,g4837);
  and AND2_322(g5498,g5449,g3460);
  and AND2_323(g1585,g1017,g1011);
  and AND2_324(g6275,g1735,g6070);
  and AND2_325(g6311,g3837,g6194);
  and AND2_326(g4671,g4645,g4641);
  and AND3_12(g4247,g1764,g4007,g1628);
  and AND2_327(g3454,g2933,g1660);
  and AND2_328(g4826,g4209,g4463);
  and AND2_329(g5162,g5088,g2105);
  and AND2_330(g5362,g4437,g5174);
  and AND2_331(g3296,g3054,g2650);
  and AND2_332(g5419,g386,g5292);
  and AND2_333(g3725,g118,g3251);
  and AND2_334(g2935,g2291,g1788);
  and AND2_335(g5452,g5315,g4612);
  and AND2_336(g6559,g1612,g6474);
  and AND2_337(g5728,g5623,g3889);
  and AND2_338(g5486,g386,g5331);
  and AND2_339(g5185,g524,g4993);
  and AND2_340(g3171,g248,g2488);
  and AND2_341(g3371,g260,g2904);
  and AND3_13(g6628,g2138,g1612,g6540);
  and AND2_342(g4165,g3927,g1352);
  and AND2_343(g4048,g414,g3388);
  and AND2_344(g4448,g3815,g4225);
  and AND2_345(g3281,g2178,g2640);
  and AND2_346(g4827,g4520,g4515);
  and AND2_347(g4333,g3964,g3284);
  and AND3_14(I2566,g749,g743,g736);
  and AND2_348(g2166,g1633,g161);
  and AND2_349(g3684,g2268,g2817);
  and AND2_350(g4396,g422,g3801);
  and AND2_351(g3338,g3162,g2914);
  and AND2_352(g2056,g1672,g1675);
  and AND2_353(g5406,g374,g5270);
  and AND2_354(g3309,g2243,g2695);
  and AND2_355(g5635,g4498,g5542);
  and AND2_356(g5682,g84,g5578);
  and AND2_357(g5487,g390,g5331);
  and AND2_358(g6123,g5702,g5958);
  and AND2_359(g6323,g3877,g6194);
  and AND2_360(g3759,g2644,g3498);
  and AND2_361(g5226,g672,g5054);
  and AND2_362(g6151,g3209,g5997);
  and AND2_363(g3449,g128,g2946);
  and AND2_364(g6648,g6579,g6234);
  and AND2_365(g5173,g512,g4993);
  and AND2_366(g5373,g161,g5250);
  and AND2_367(g4181,g3939,g1381);
  and AND2_368(g2720,g2422,g1919);
  and AND2_369(g4685,g4591,g2079);
  and AND2_370(g5169,g5093,g1375);
  and AND2_371(g5369,g143,g5247);
  and AND2_372(g5602,g594,g5515);
  and AND4_3(g2834,g1263,g1257,g1270,I4040);
  and AND2_373(g3362,g3031,g2740);
  and AND2_374(g6343,g6268,g6078);
  and AND2_375(g2121,g1632,g754);
  and AND2_376(g2670,g2029,g1503);
  and AND2_377(g6693,g6618,g6617);
  and AND2_378(g1633,g716,g152);
  and AND2_379(g6334,g3858,g6212);
  and AND2_380(g3728,g326,g3441);
  and AND2_381(g6555,g1838,g6469);
  and AND2_382(g3730,g328,g3441);
  and AND2_383(g2909,g606,g2092);
  and AND2_384(g4041,g461,g3388);
  and AND2_385(g3425,g2296,g3208);
  and AND2_386(g6313,g3841,g6194);
  and AND2_387(g5940,g5115,g5794);
  and AND2_388(g4673,g4656,g4654);
  and AND2_389(g5188,g1043,g4894);
  and AND2_390(g6908,g6907,g3886);
  and AND2_391(g5216,g563,g5025);
  and AND2_392(g6094,g1177,g5753);
  and AND2_393(g4168,g3925,g1355);
  and AND2_394(g4368,g3998,g3363);
  and AND2_395(g5671,g54,g5572);
  and AND2_396(g3678,g2256,g2802);
  and AND2_397(g5428,g394,g5300);
  and AND2_398(g4058,g3424,g1246);
  and AND2_399(g3635,g2473,g3079);
  and AND2_400(g2860,g710,g2296);
  and AND2_401(g3682,g2772,g2430);
  and AND2_402(g3305,g2960,g2296);
  and AND2_403(g5910,g5816,g5667);
  and AND2_404(g3755,g2604,g3481);
  and AND2_405(g2659,g1686,g2296);
  and AND2_406(g5883,g5824,g3752);
  and AND2_407(g3373,g3118,g2927);
  and AND2_408(g5217,g4866,g5092);
  and AND2_409(g4863,g4777,g2874);
  and AND2_410(g3283,g2609,g2622);
  and AND2_411(g3602,g2688,g2663);
  and AND3_15(I2574,g804,g798,g791);
  and AND2_412(g5165,g508,g4993);
  and AND2_413(g6777,g6762,g3488);
  and AND3_16(g3718,g1743,g3140,g1157);
  and AND2_414(g3767,g2706,g3504);
  and AND2_415(g4688,g1474,g4568);
  and AND2_416(g1784,g858,g889);
  and AND2_417(g2853,g836,g2021);
  and AND2_418(g6799,g4948,g6782);
  and AND2_419(g2794,g2544,g1994);
  and AND2_420(g3203,g2497,g2565);
  and AND2_421(g6132,g3752,g5880);
  and AND2_422(g6238,g528,g5886);
  and AND2_423(g6153,g3216,g5997);
  and AND2_424(g4183,g3965,g1391);
  and AND2_425(g4383,g453,g3796);
  and AND2_426(g6558,g1842,g6474);
  and AND2_427(g5181,g449,g4877);
  and AND2_428(g3689,g3162,g2826);
  and AND2_429(g4588,g2419,g4273);
  and AND2_430(g5197,g465,g4967);
  and AND2_431(g4161,g3931,g2087);
  and AND2_432(g4361,g3995,g3354);
  and AND2_433(g3671,g2760,g2405);
  and AND2_434(g4051,g449,g3388);
  and AND2_435(g6092,g1123,g5731);
  and AND2_436(g4346,g157,g3773);
  and AND2_437(g2323,g471,g1358);
  and AND2_438(g5562,g5228,g5457);
  and AND2_439(g3910,g3546,g1049);
  and AND2_440(g3609,g2706,g2678);
  and AND2_441(g6262,g516,g5901);
  and AND3_17(g6736,g6712,g754,g5237);
  and AND2_442(g3758,g545,g3461);
  and AND2_443(g4043,g457,g3388);
  and AND2_444(g3365,g254,g2892);
  and AND3_18(g5441,g4537,g5251,g1558);
  and AND2_445(g5673,g59,g5573);
  and AND2_446(g4347,g3986,g3320);
  and AND2_447(g3133,g236,g2410);
  and AND2_448(g3333,g2264,g2728);
  and AND2_449(g3774,g3016,g3510);
  and AND2_450(g4697,g4589,g1363);
  and AND2_451(g3780,g3043,g3519);
  and AND3_19(g6737,g6714,g760,g5237);
  and AND2_452(g6077,g5824,g1735);
  and AND2_453(g3662,g2544,g3114);
  and AND2_454(g6643,g6574,g6229);
  and AND2_455(g3290,g2213,g2664);
  and AND2_456(g6634,g1595,g6545);
  and AND2_457(g3816,g3434,g861);
  and AND2_458(g2113,g1576,g1535);
  and AND2_459(g6099,g1222,g5753);
  and AND2_460(g6304,g5915,g6165);
  and AND2_461(g3181,g254,g2509);
  and AND2_462(g3381,g3128,g1998);
  and AND2_463(g3685,g2256,g2818);
  and AND2_464(g3700,g2276,g2837);
  and AND2_465(g3421,g622,g2846);
  and AND2_466(g5569,g5348,g3772);
  and AND2_467(g4460,g4218,g1539);
  and AND2_468(g4597,g3694,g4286);
  and AND2_469(g6613,g932,g6554);
  and AND2_470(g4739,g2850,g4579);
  and AND2_471(g6269,g524,g5908);
  and AND2_472(g4937,g166,g4732);
  and AND2_473(g4668,g4642,g4638);
  and AND2_474(g3631,g2631,g2324);
  and AND2_475(g2160,g1624,g929);
  and AND2_476(g4390,g418,g3799);
  and AND2_477(g3301,g218,g2866);
  and AND2_478(g4501,g4250,g1671);
  and AND2_479(g4156,g3926,g2078);
  and AND2_480(g4356,g175,g3779);
  and AND2_481(g4942,g175,g4736);
  and AND2_482(g5183,g418,g4950);
  and AND2_483(g4163,g374,g3892);
  and AND2_484(g5023,g3935,g4804);
  and AND2_485(g4363,g402,g3786);
  and AND2_486(g4032,g441,g3388);
  and AND2_487(g4053,g3387,g1415);
  and AND2_488(g4453,g4238,g1858);
  and AND2_489(g5161,g5095,g4535);
  and AND2_490(g3669,g2234,g2790);
  and AND2_491(g5361,g4435,g5168);
  and AND2_492(g3368,g2822,g2923);
  and AND2_493(g6135,g5584,g5958);
  and AND2_494(g5665,g361,g5570);
  and AND2_495(g6831,g6812,g5975);
  and AND2_496(g5451,g5251,g4544);
  and AND2_497(g6288,g5615,g6160);
  and AND2_498(g4157,g3830,g1533);
  and AND2_499(g4357,g3990,g3342);
  and AND2_500(g5146,g184,g5099);
  and AND2_501(g6916,g6903,g6901);
  and AND2_502(g5633,g4496,g5539);
  and AND2_503(g3505,g2924,g1749);
  and AND2_504(g6749,g6735,g6734);
  and AND2_505(g6798,g4946,g6781);
  and AND2_506(g5944,g5778,g5403);
  and AND2_507(g5240,g293,g4915);
  and AND2_508(g5043,g3941,g4805);
  and AND3_20(g5443,g4537,g5251,g2307);
  and AND2_509(g6302,g5740,g6164);
  and AND2_510(g6719,g4518,g6665);
  and AND2_511(g2092,g642,g1570);
  and AND2_512(g4683,g4585,g2066);
  and AND2_513(g5681,g79,g5577);
  and AND2_514(g3688,g2783,g2457);
  and AND2_515(g4735,g2018,g4577);
  and AND2_516(g6265,g520,g5903);
  and AND2_517(g4782,g1624,g4623);
  and AND2_518(g4661,g4637,g4634);
  and AND2_519(g4949,g193,g4753);
  and AND2_520(g3326,g2734,g1891);
  and AND2_521(g6770,g6754,g3482);
  and AND2_522(g3760,g548,g3465);
  and AND2_523(g5936,g5113,g5788);
  and AND2_524(g4039,g402,g3388);
  and AND2_525(g5317,g148,g4869);
  and AND2_526(g3383,g3128,g2004);
  and AND2_527(g5601,g5052,g5518);
  and AND2_528(g3608,g2599,g2308);
  and AND2_529(g3924,g3505,g471);
  and AND2_530(g4583,g1808,g4267);
  and AND2_531(g3161,g2397,g2470);
  and AND2_532(g2339,g1603,g197);
  and AND2_533(g3361,g3150,g1950);
  and AND2_534(g4616,g4231,g3761);
  and AND2_535(g3665,g2748,g2378);
  and AND2_536(g3127,g224,g2394);
  and AND2_537(g3327,g2772,g2906);
  and AND2_538(g3146,g2370,g2446);
  and AND2_539(g3633,g2497,g3076);
  and AND2_540(g5937,g5775,g5392);
  and AND2_541(g3103,g212,g2353);
  and AND2_542(g3303,g2722,g2890);
  and AND2_543(g5668,g49,g5571);
  and AND2_544(g6338,g6251,g6067);
  and AND2_545(g5190,g426,g4950);
  and AND2_546(g5501,g5454,g3478);
  and AND2_547(g2551,g715,g1826);
  and AND2_548(g5156,g434,g4877);
  and AND2_549(g5356,g5265,g1902);
  and AND2_550(g4277,g3936,g942);
  and AND2_551(g5942,g5117,g5797);
  and AND2_552(g4789,g3551,g4632);
  and AND2_553(g3316,g2748,g2894);
  and AND2_554(g3434,g2850,g857);
  and AND2_555(g5954,g5121,g5813);
  and AND2_556(g5163,g402,g4950);
  and AND2_557(g6098,g1209,g5753);
  and AND2_558(g3147,g2419,g59);
  and AND2_559(g5363,g4439,g5179);
  and AND2_560(g3681,g2234,g2806);
  and AND2_561(g5053,g4599,g4808);
  and AND2_562(g3697,g2796,g2481);
  and AND2_563(g5157,g496,g4904);
  and AND2_564(g5357,g398,g5220);
  and AND3_21(g4244,g1749,g4004,g1609);
  and AND2_565(g4340,g3972,g3291);
  and AND2_566(g3936,g3551,g940);
  and AND2_567(g3117,g218,g2367);
  and AND2_568(g3317,g2722,g2895);
  and AND2_569(g4035,g437,g3388);
  and AND2_570(g918,g610,g602);
  and AND2_571(g6086,g1143,g5742);
  and AND2_572(g4214,g1822,g4045);
  and AND2_573(g1620,g1056,g1084);
  and AND2_574(g3784,g114,g3251);
  and AND2_575(g2916,g1030,g2113);
  and AND2_576(g3479,g345,g2957);
  and AND2_577(g6131,g5593,g5975);
  and AND2_578(g3668,g2568,g3124);
  and AND2_579(g6331,g3891,g6212);
  and AND2_580(g4236,g654,g3907);
  and AND2_581(g3294,g139,g2870);
  and AND2_582(g5949,g5119,g5805);
  and AND2_583(g3190,g260,g2535);
  and AND2_584(g6766,g6750,g2986);
  and AND2_585(g3156,g242,g2464);
  and AND2_586(g3356,g248,g2888);
  and AND2_587(g5646,g4502,g5544);
  and AND2_588(g2873,g1845,g1861);
  and AND2_589(g6748,g6733,g6732);
  and AND2_590(g5603,g5504,g4911);
  and AND2_591(g5484,g378,g5331);
  and AND2_592(g4928,g148,g4723);
  and AND2_593(g3704,g2276,g2841);
  and AND2_594(g4464,g4272,g1937);
  and AND2_595(g4785,g2160,g4625);
  and AND2_596(g6091,g1161,g5753);
  and AND2_597(g3810,g625,g3421);
  and AND2_598(g5952,g5120,g5809);
  and AND2_599(g5616,g5505,g4929);
  and AND2_600(g6718,g4511,g6661);
  and AND2_601(g6767,g6754,g2986);
  and AND2_602(g3157,g2422,g2467);
  and AND2_603(g3357,g242,g2889);
  and AND2_604(g4489,g2166,g4206);
  and AND2_605(g2770,g2518,g1972);
  and AND2_606(g4471,g4253,g332);
  and AND2_607(g5503,g366,g5384);
  and AND2_608(g3626,g3031,g2727);
  and AND2_609(g4038,g430,g3388);
  and AND2_610(g5617,g5061,g5524);
  and AND2_611(g3683,g3150,g2813);
  and AND2_612(g4836,g4527,g4523);
  and AND2_613(g2138,g1639,g809);
  and AND2_614(g3661,g2234,g2778);
  and AND2_615(g6247,g504,g5893);
  and AND2_616(g3627,g2473,g3067);
  and AND2_617(g5945,g5118,g5801);
  and AND2_618(g2808,g2009,g1581);
  and AND2_619(g3292,g2214,g2667);
  and AND2_620(g3646,g2179,g2756);
  and AND2_621(g2759,g2473,g1966);
  and AND2_622(g6910,g6892,g6891);
  and AND2_623(g3603,g2370,g3019);
  and AND2_624(g3484,g349,g2958);
  and AND2_625(g5482,g370,g5331);
  and AND2_626(g3702,g2284,g2839);
  and AND2_627(g6066,g5824,g1721);
  and AND2_628(g5214,g562,g5025);
  and AND2_629(g3616,g2397,g3049);
  and AND2_630(g6055,g5824,g1696);
  and AND2_631(g6133,g5723,g5975);
  and AND2_632(g5663,g4513,g5550);
  and AND2_633(g6333,g3896,g6212);
  and AND2_634(g2419,g1808,g54);
  and AND2_635(g3764,g551,g3480);
  and AND2_636(g5402,g370,g5266);
  and AND2_637(g5236,g269,g4915);
  and AND2_638(g4708,g578,g4541);
  and AND2_639(g5556,g5015,g5445);
  and AND2_640(g4219,g3911,g1655);
  and AND2_641(g3277,g2174,g2625);
  and AND2_642(g3617,g2609,g2317);
  and AND2_643(g6093,g1177,g5742);
  and AND2_644(g2897,g1030,g2062);
  and AND2_645(g6256,g1696,g6040);
  and AND2_646(g4176,g386,g3901);
  and AND2_647(g6816,g6784,g3346);
  and AND2_648(g4829,g4526,g4522);
  and AND2_649(g6263,g1711,g6052);
  and AND2_650(g5194,g586,g4874);
  and AND2_651(g3709,g2284,g2845);
  and AND2_652(g5557,g5016,g5448);
  and AND2_653(g3340,g2772,g2915);
  and AND2_654(g6631,g1838,g6545);
  and AND2_655(g3907,g650,g3522);
  and AND2_656(g4177,g3933,g1372);
  and AND2_657(g5948,g5779,g5407);
  and AND2_658(g4377,g457,g3791);
  and AND2_659(g3690,g2276,g2827);
  and AND2_660(g5955,g5782,g5420);
  and AND2_661(g5350,g5325,g3453);
  and AND2_662(g4199,g628,g3810);
  and AND2_663(g5438,g5224,g3769);
  and AND2_664(g2868,g1316,g1861);
  and AND2_665(g3310,g224,g2871);
  and AND2_666(g4797,g4593,g4643);
  and AND2_667(g5212,g561,g5025);
  and AND2_668(g3663,g2215,g2779);
  and AND2_669(g2793,g2568,g1991);
  and AND2_670(g2015,g616,g1419);
  and AND2_671(g4344,g3981,g3306);
  and AND2_672(g5229,g545,g4980);
  and AND2_673(g6772,g6746,g3312);
  and AND2_674(g3762,g2672,g3500);
  and AND2_675(g4694,g1481,g4578);
  and AND2_676(g3657,g2734,g2357);
  and AND2_677(g2721,g2397,g1922);
  and AND2_678(g4488,g1633,g4202);
  and AND2_679(g4701,g4596,g1378);
  and AND2_680(g3928,g3512,g478);
  and AND3_22(g6474,g2138,g2036,g6397);
  and AND2_681(g3899,g323,g3441);
  and AND2_682(g3464,g341,g2956);
  and AND2_683(g5620,g5507,g4938);
  and AND2_684(g4870,g4779,g1884);
  and AND2_685(g3295,g2660,g2647);
  and AND2_686(g2671,g2263,g2296);
  and AND2_687(g1576,g1101,g1094);
  and AND2_688(g3844,g3540,g1665);
  and AND3_23(g1716,g821,g774,g784);
  and AND2_689(g3089,g212,g2336);
  and AND2_690(g3731,g331,g3441);
  and AND2_691(g3489,g2607,g1861);
  and AND2_692(g5192,g1046,g4894);
  and AND2_693(g5485,g382,g5331);
  and AND2_694(g5941,g5777,g5399);
  and AND2_695(g4230,g3756,g1861);
  and AND2_696(g6126,g5711,g5958);
  and AND2_697(g6326,g3833,g6194);
  and AND2_698(g4033,g426,g3388);
  and AND2_699(g3814,g913,g3546);
  and AND2_700(g2758,g2497,g1963);
  and AND2_701(g3350,g3150,g1928);
  and AND2_702(g2861,g2120,g1654);
  and AND2_703(g6924,g6920,g6919);
  and AND2_704(g5176,g410,g4950);
  and AND2_705(g4395,g445,g3800);
  and AND2_706(g5376,g170,g5255);
  and AND2_707(g5911,g5817,g5670);
  and AND2_708(g2846,g619,g2015);
  and AND2_709(g6127,g5714,g5975);
  and AND2_710(g6327,g3884,g6212);
  and AND2_711(g5225,g669,g5054);
  and AND2_712(g4342,g3978,g3299);
  and AND2_713(g6146,g3192,g5997);
  and AND2_714(g6346,g6274,g6087);
  and AND2_715(g2018,g1423,g1254);
  and AND2_716(g4354,g437,g3777);
  and AND4_4(I5352,g3529,g3531,g3535,g3538);
  and AND2_717(g5177,g445,g4877);
  and AND2_718(g6240,g4205,g5888);
  and AND2_719(g3620,g2422,g3060);
  and AND2_720(g1027,g598,g567);
  and AND2_721(g2685,g2370,g1887);
  and AND2_722(g2700,g2370,g1908);
  and AND2_723(g2021,g835,g1436);
  and AND2_724(g6316,g3855,g6194);
  and AND2_725(g5898,g5800,g5647);
  and AND2_726(g4401,g426,g3802);
  and AND2_727(g1514,g1017,g1011);
  and AND2_728(g5900,g5804,g5658);
  and AND2_729(g2950,g2156,g1612);
  and AND2_730(g4761,g4567,g1674);
  and AND2_731(g5245,g297,g4915);
  and AND2_732(g1763,g478,g1119);
  and AND2_733(g4828,g4510,g4508);
  and AND2_734(g3298,g2231,g2679);
  and AND2_735(g4830,g4529,g4525);
  and AND2_736(g5144,g166,g5099);
  and AND2_737(g4592,g3147,g4281);
  and AND2_738(g6914,g6895,g6893);
  and AND2_739(g2101,g1001,g1543);
  and AND2_740(g5488,g394,g5331);
  and AND2_741(g4932,g157,g4727);
  and AND2_742(g1416,g913,g266);
  and AND2_743(g5701,g5683,g3813);
  and AND2_744(g6317,g3862,g6194);
  and AND2_745(g5215,g4864,g5090);
  and AND2_746(g5951,g5780,g5411);
  and AND2_747(g4677,g4652,g4646);
  and AND2_748(g3176,g2422,g2494);
  and AND2_749(g3376,g3104,g1979);
  and AND2_750(g3286,g2196,g2656);
  and AND2_751(g3765,g554,g3485);
  and AND2_752(g4349,g441,g3775);
  and AND2_753(g6060,g5824,g1703);
  and AND4_5(g1595,g729,g719,g766,I2566);
  and AND4_6(I5359,g3518,g3521,g3526,g3530);
  and AND2_754(g3610,g2397,g3034);
  and AND3_24(g6739,g6715,g815,g5242);
  and AND4_7(g1612,g784,g774,g821,I2574);
  and AND2_755(g3324,g230,g2875);
  and AND2_756(g6079,g1236,g5753);
  and AND2_757(g5122,g193,g4662);
  and AND2_758(g3377,g3118,g2931);
  and AND2_759(g4352,g3988,g3331);
  and AND2_760(g4867,g4811,g3872);
  and AND2_761(g6156,g2591,g6015);
  and AND2_762(g3287,g135,g2865);
  and AND2_763(g5096,g4794,g4647);
  and AND2_764(g4186,g3973,g1395);
  and AND2_765(g5496,g5446,g3457);
  and AND2_766(g6250,g1692,g6036);
  and AND2_767(g4170,g382,g3900);
  and AND3_25(g4280,g2138,g1764,g4007);
  and AND2_768(g3144,g236,g2440);
  and AND2_769(g3344,g242,g2885);
  and AND2_770(g5142,g148,g5099);
  and AND2_771(g3819,g964,g3437);
  and AND2_772(g6912,g6899,g6897);
  and AND2_773(g3694,g3147,g64);
  and AND2_774(g6157,g3158,g5997);
  and AND2_775(g5481,g366,g5331);
  and AND2_776(g3701,g2268,g2838);
  and AND2_777(g5497,g5447,g3458);
  and AND2_778(g5154,g500,g4993);
  and AND2_779(g5354,g5249,g2903);
  and AND2_780(g4461,g4241,g2919);
  and AND2_781(g4756,g3816,g4587);
  and AND2_782(g4046,I5351,I5352);
  and AND2_783(g5218,g564,g5025);
  and AND2_784(g3650,g2660,g2347);
  and AND2_785(g4345,g3982,g3308);
  and AND2_786(g3336,g2760,g1911);
  and AND2_787(g3768,g3448,g1528);
  and AND2_788(g4159,g370,g3890);
  and AND2_789(g4359,g434,g3782);
  and AND2_790(g3806,g3384,g2024);
  and AND2_791(g4416,g3905,g1481);
  and AND2_792(g3887,g3276,g1861);
  and AND2_793(g3122,g2435,g1394);
  and AND2_794(g2732,g2449,g1940);
  and AND2_795(g4047,g453,g3388);
  and AND2_796(g6646,g6577,g6232);
  and AND3_26(g3433,g1359,g2831,g905);
  and AND2_797(g5953,g5781,g5415);
  and AND2_798(g6084,g1123,g5753);
  and AND2_799(g6603,g6581,g6236);
  and AND2_800(g4874,g582,g4708);
  and AND2_801(g5677,g69,g5575);
  and AND2_802(g3195,g2473,g2541);
  and AND2_803(g3337,g2796,g2913);
  and AND3_27(I4040,g1279,g2025,g1267);
  and AND2_804(g5149,g4910,g1480);
  and AND2_805(g5349,g5324,g3451);
  and AND2_806(g5198,g558,g5025);
  and AND2_807(g5398,g366,g5261);
  and AND2_808(g1570,g634,g1027);
  and AND2_809(g6647,g6578,g6233);
  and AND2_810(g1691,g821,g774);
  and AND2_811(g3692,g2268,g2829);
  and AND2_812(g3726,g119,g3251);
  and AND2_813(g3154,g2039,g1410);
  and AND2_814(g4800,g4648,g4296);
  and AND2_815(g5152,g430,g4950);
  and AND2_816(g6320,g3869,g6194);
  and AND2_817(g5211,g4860,g5086);
  and AND2_818(g5186,g422,g4950);
  and AND2_819(g5599,g5049,g5512);
  and AND2_820(g4490,g2941,g4210);
  and AND2_821(g3293,g212,g2864);
  and AND2_822(g6771,g6758,g3483);
  and AND2_823(g3329,g2748,g2907);
  and AND2_824(g5170,g5091,g2111);
  and AND2_825(g4456,g3829,g4229);
  and AND2_826(g6299,g5530,g6163);
  and AND2_827(g4348,g3987,g3322);
  and AND2_828(g3727,g122,g3251);
  and AND2_829(g2937,g2160,g931);
  and AND2_830(g4355,g430,g3778);
  and AND2_831(g5939,g5776,g5395);
  and AND3_28(g2294,g1716,g791,g798);
  and AND2_832(g4698,g4586,g2106);
  and AND2_833(g5483,g374,g5331);
  and AND2_834(g3703,g2284,g2840);
  and AND3_29(g6738,g6713,g809,g5242);
  and AND2_835(g2156,g815,g1642);
  and AND2_836(g6244,g4759,g5891);
  and AND2_837(g2356,g1603,g269);
  and AND2_838(g6140,g5587,g5975);
  and AND2_839(g3953,g3554,g188);
  and AND2_840(g6340,g6257,g6069);
  and AND2_841(g5187,g457,g4877);
  and AND2_842(g1628,g815,g809);
  and AND2_843(g4167,g378,g3898);
  and AND2_844(g6082,g1123,g5742);
  and AND2_845(g4367,g193,g3788);
  and AND2_846(g4872,g4760,g1549);
  and AND2_847(g4057,g422,g3388);
  and AND2_848(g5904,g5812,g5664);
  and AND2_849(g5200,g559,g5025);
  and AND2_850(g4457,g4261,g2902);
  and AND2_851(g5446,g4537,g5241);
  and AND2_852(g3349,g2783,g1925);
  and AND2_853(g2053,g1094,g1675);
  and AND2_854(g5145,g175,g5099);
  and AND2_855(g6915,g6906,g6905);
  and AND2_856(g4834,g4534,g4531);
  and AND2_857(g4686,g4590,g1348);
  and AND2_858(g5191,g461,g4877);
  and AND2_859(g3699,g2276,g2836);
  and AND2_860(g4598,g1978,g4253);
  and AND2_861(g5637,g4499,g5543);
  and AND2_862(g5159,g536,g4967);
  and AND2_863(g5359,g4428,g5155);
  and AND2_864(g4253,g1861,g3819);
  and AND2_865(g3644,g2197,g2755);
  and AND2_866(g3319,g2688,g2675);
  and AND2_867(g3352,g2796,g2920);
  and AND2_868(g5047,g3954,g4806);
  and AND3_30(g5447,g4545,g5256,g2311);
  and AND2_869(g4687,g4493,g1542);
  and AND2_870(g3186,g2449,g2515);
  and AND2_871(g3170,g254,g2485);
  and AND2_872(g3614,g2998,g2691);
  and AND2_873(g3325,g224,g2876);
  and AND2_874(g4341,g3977,g3297);
  and AND2_875(g2782,g2518,g1985);
  and AND2_876(g6295,g5379,g6162);
  and AND2_877(g3280,g2177,g2637);
  and AND2_878(g5017,g4784,g1679);
  and AND2_879(g4691,g4581,g2098);
  and AND2_880(g5935,g5112,g5784);
  and AND2_881(g2949,g830,g1861);
  and AND4_8(I5351,g3511,g3517,g3520,g3525);
  and AND2_882(g5234,g197,g4915);
  and AND2_883(g3636,g2701,g2327);
  and AND3_31(g2292,g1706,g736,g743);
  and AND2_884(g6089,g1143,g5731);
  and AND2_885(g6731,g6717,g4427);
  and AND2_886(g6557,g1595,g6469);
  and AND2_887(g4358,g3991,g3343);
  and AND2_888(g2084,g1577,g1563);
  and AND2_889(g2850,g2018,g1255);
  and AND2_890(g5213,g4862,g5087);
  and AND2_891(g6254,g532,g5897);
  and AND2_892(g6150,g3204,g6015);
  and AND2_893(g5902,g5808,g5661);
  and AND2_894(g3145,g2397,g2443);
  and AND2_895(g3345,g236,g2886);
  and AND2_896(g6773,g6762,g2986);
  and AND2_897(g3763,g3064,g3501);
  and AND2_898(g3191,g2497,g2538);
  and AND2_899(g4180,g3929,g2119);
  and AND2_900(g5166,g541,g4967);
  and AND2_901(g3637,g2822,g2752);
  and AND2_902(g4832,g4517,g4512);
  and AND2_903(g6769,g6758,g2986);
  and AND2_904(g3307,g2242,g2692);
  and AND2_905(g3359,g2822,g2922);
  and AND2_906(g4794,g4593,g949);
  and AND2_907(g3757,g2619,g3487);
  and AND2_908(g3522,g646,g2909);
  and AND2_909(g3315,g2701,g1875);
  and AND2_910(g3642,g3054,g2754);
  and AND2_911(g3654,g2518,g3100);
  and AND2_912(g5619,g5064,g5527);
  and AND2_913(g5167,g5011,g1556);
  or OR2_0(g3880,g3658,g3665);
  or OR2_1(g4440,g4371,g4038);
  or OR2_2(g3978,g3655,g3117);
  or OR2_3(g6788,g3760,g6767);
  or OR2_4(g3935,g3464,g2868);
  or OR2_5(g3982,g3663,g3127);
  or OR4_0(I8376,g6315,g6126,g6129,g6146);
  or OR2_6(g5625,g5495,g3281);
  or OR2_7(g6298,g6255,g6093);
  or OR3_0(g6485,I8393,I8394,I8395);
  or OR2_8(g4655,g4368,g3660);
  or OR2_9(g6252,g5905,g2381);
  or OR2_10(g6176,g6068,g6033);
  or OR4_1(I8377,g6150,g6324,g5180,g5181);
  or OR2_11(g6286,g6238,g6079);
  or OR2_12(g3851,g3681,g3146);
  or OR2_13(g3964,g3634,g3089);
  or OR2_14(g5659,g5551,g5398);
  or OR2_15(g2928,g2100,g1582);
  or OR2_16(g6287,g6241,g6082);
  or OR2_17(g3989,g3679,g3144);
  or OR2_18(g5374,g5215,g4947);
  or OR2_19(g3971,g3644,g3099);
  or OR2_20(g6781,g6718,g6748);
  or OR2_21(g3598,g2808,g2821);
  or OR2_22(g4641,g4347,g3627);
  or OR2_23(g4450,g4389,g4047);
  or OR2_24(g3740,g3335,g2747);
  or OR4_2(I8136,g6015,g6212,g4950,g4877);
  or OR2_25(g5628,g5498,g3292);
  or OR2_26(g5630,g5501,g3309);
  or OR2_27(g6114,g5904,g5604);
  or OR2_28(g5323,g5098,g4802);
  or OR2_29(g5666,g5555,g5406);
  or OR4_3(I8137,g4894,g4904,g4993,g4967);
  or OR3_1(I8395,g5182,g5200,g6280);
  or OR2_30(g3879,g3704,g3195);
  or OR4_4(I9057,g6320,g6828,g6830,g6153);
  or OR2_31(g4092,g3311,g2721);
  or OR4_5(I8081,g4894,g4904,g4993,g4967);
  or OR2_32(g4864,g4744,g4490);
  or OR3_2(g6845,I9064,I9065,I9066);
  or OR2_33(g5372,g5213,g4942);
  or OR2_34(g5693,g5632,g5481);
  or OR2_35(g5804,g5371,g5603);
  or OR2_36(g6142,g5909,g3806);
  or OR2_37(I8129,g4915,g5025);
  or OR4_6(g6481,I8367,I8368,I8369,I8370);
  or OR2_38(g4651,g4357,g3643);
  or OR2_39(g4285,g3490,g3887);
  or OR2_40(g4500,g4243,g2010);
  or OR3_3(g5202,g4904,g4914,g4894);
  or OR2_41(g3750,g3372,g2794);
  or OR2_42(g6267,g2953,g5884);
  or OR2_43(g4231,g3997,g4000);
  or OR2_44(g6676,g6631,g6555);
  or OR2_45(g6293,g6244,g6085);
  or OR2_46(g4205,g3843,g541);
  or OR2_47(g4634,g4341,g3615);
  or OR4_7(I8349,I8345,I8346,I8347,I8348);
  or OR2_48(g6703,g6692,g4831);
  or OR2_49(g3884,g3666,g3671);
  or OR2_50(g4444,g4378,g4042);
  or OR2_51(g4862,g4739,g4489);
  or OR4_8(I8119,g5202,g4993,g4967,g4980);
  or OR2_52(g3988,g3678,g3143);
  or OR2_53(g5674,g5558,g5419);
  or OR2_54(g6747,g6614,g6731);
  or OR2_55(g6855,g6851,g2085);
  or OR2_56(I8211,g4915,g5025);
  or OR4_9(I8386,g6152,g6327,g5183,g5177);
  or OR2_57(g5680,g5562,g5429);
  or OR2_58(g4946,g4830,g4833);
  or OR2_59(I8370,g5214,g6358);
  or OR2_60(g4436,g4359,g4035);
  or OR3_4(I8387,g5178,g5209,g6281);
  or OR2_61(g6274,g5682,g5956);
  or OR2_62(g6426,g6288,g6119);
  or OR2_63(g6170,g6061,g6014);
  or OR2_64(g3996,g3691,g3171);
  or OR4_10(I8345,g6326,g6135,g6140,g6157);
  or OR2_65(g5623,g5503,g5357);
  or OR3_5(g6483,I8385,I8386,I8387);
  or OR2_66(g4653,g4361,g3652);
  or OR2_67(g3878,g3703,g3191);
  or OR2_68(g6790,g3765,g6773);
  or OR4_11(I8359,g5232,g5236,g5216,g5226);
  or OR2_69(g4752,g4452,g4155);
  or OR2_70(g6461,g6353,g6351);
  or OR2_71(g3981,g3661,g3123);
  or OR2_72(g5024,g4793,g4600);
  or OR2_73(g4233,g3912,g471);
  or OR2_74(g4454,g4395,g4051);
  or OR2_75(g5672,g5557,g5414);
  or OR2_76(g5077,g1612,g4694);
  or OR2_77(g5231,g5048,g672);
  or OR2_78(g6307,g6262,g6096);
  or OR2_79(g3744,g3345,g2759);
  or OR2_80(g6251,g5668,g5939);
  or OR2_81(g6447,g6340,g5938);
  or OR4_12(I8128,g5202,g4993,g4967,g4980);
  or OR2_82(g3864,g3693,g3176);
  or OR2_83(g5044,g4797,g4602);
  or OR2_84(g4745,g4468,g4569);
  or OR2_85(g6272,g5679,g5953);
  or OR2_86(g5014,g4785,g4583);
  or OR2_87(g3871,g3701,g3186);
  or OR4_13(I7970,g6015,g6212,g4950,g4877);
  or OR4_14(I8348,g5229,g5234,g5218,g5225);
  or OR2_88(g6554,g6337,g6466);
  or OR4_15(I7987,g6194,g5958,g5975,g5997);
  or OR2_89(g5916,g5728,g3781);
  or OR4_16(I8118,g6015,g6212,g4950,g4877);
  or OR4_17(I8367,g6313,g6124,g6127,g6144);
  or OR2_90(g6456,g6346,g5954);
  or OR4_18(I8393,g6317,g6130,g6133,g6151);
  or OR2_91(g4086,g3310,g2720);
  or OR2_92(g1589,g1059,g1045);
  or OR2_93(g6118,g5911,g5619);
  or OR2_94(g6167,g6056,g6039);
  or OR2_95(g3862,g3632,g3641);
  or OR2_96(g6457,g6352,g6347);
  or OR2_97(g4635,g4342,g3616);
  or OR2_98(g6549,g6473,g4247);
  or OR2_99(g6686,g6259,g6645);
  or OR2_100(g5532,g5350,g3278);
  or OR4_19(g6670,g6557,g6634,g4410,g2948);
  or OR2_101(g5012,g4782,g4580);
  or OR2_102(g4059,g3466,g3425);
  or OR2_103(g5281,g5074,g5124);
  or OR4_20(I8358,g5192,g5153,g5158,g5197);
  or OR2_104(g6687,g6260,g6646);
  or OR2_105(g3749,g3371,g2793);
  or OR2_106(g5808,g5373,g5616);
  or OR2_107(g6691,g6275,g6603);
  or OR2_108(g3873,g3649,g3657);
  or OR2_109(g3869,g3642,g3650);
  or OR2_110(g6659,g6634,g6631);
  or OR2_111(g4430,g4349,g4015);
  or OR2_112(g6239,g2339,g6073);
  or OR2_113(g6545,g6468,g4244);
  or OR2_114(g4638,g4345,g3620);
  or OR2_115(g6794,g6777,g3333);
  or OR2_116(g6931,g6741,g6929);
  or OR2_117(g3990,g3684,g3155);
  or OR2_118(g5385,g3992,g5318);
  or OR2_119(g3888,g3672,g3682);
  or OR2_120(g5470,g5359,g5142);
  or OR2_121(g6300,g6253,g6091);
  or OR2_122(g4455,g4396,g4052);
  or OR3_6(g6750,g6670,g6625,g6736);
  or OR2_123(g5678,g5560,g5428);
  or OR2_124(g3745,g3356,g2770);
  or OR2_125(g6440,g6336,g5935);
  or OR2_126(g3865,g3637,g3648);
  or OR2_127(g3833,g3602,g3608);
  or OR2_128(g4021,g3558,g2949);
  or OR2_129(g3896,g3689,g3697);
  or OR2_130(g5535,g5353,g3300);
  or OR2_131(g5015,g4787,g4588);
  or OR2_132(g4631,g4340,g3611);
  or OR2_133(g5246,g5077,g2080);
  or OR2_134(g6792,g6770,g3321);
  or OR4_21(I7980,g5202,g4993,g4967,g4980);
  or OR4_22(I8360,I8356,I8357,I8358,I8359);
  or OR2_135(g4441,g4372,g4039);
  or OR2_136(g6113,g5902,g5601);
  or OR3_7(g5388,g5318,g1589,g3491);
  or OR2_137(I8379,g5212,g6357);
  or OR2_138(g5430,g5161,g4873);
  or OR2_139(g4458,g4401,g4057);
  or OR2_140(g3748,g3366,g2782);
  or OR2_141(g6264,g5675,g5948);
  or OR2_142(g4074,g3301,g2699);
  or OR2_143(g6450,g6341,g5940);
  or OR2_144(g4080,g3302,g2700);
  or OR2_145(g5066,g4668,g4672);
  or OR2_146(g6179,g6077,g6051);
  or OR4_23(I8209,g6015,g6212,g4950,g4877);
  or OR2_147(g6289,g6240,g6081);
  or OR2_148(g6658,g6132,g6620);
  or OR2_149(g6271,g2955,g5885);
  or OR2_150(g5662,g5553,g5402);
  or OR2_151(g5018,g4791,g4597);
  or OR2_152(I7972,g4915,g5025);
  or OR3_8(g5467,g3868,g5318,g3992);
  or OR2_153(g5816,g5378,g5620);
  or OR2_154(g5700,g5663,g5488);
  or OR2_155(g4451,g4390,g4048);
  or OR2_156(g6864,g6852,g2089);
  or OR2_157(g5817,g5380,g5621);
  or OR2_158(g3883,g3709,g3203);
  or OR2_159(g5605,g3575,g5500);
  or OR3_9(I9059,g5185,g5198,g6279);
  or OR2_160(g4443,g4377,g4041);
  or OR2_161(g4434,g4355,g4033);
  or OR2_162(g5669,g5556,g5410);
  or OR2_163(g5368,g5201,g4932);
  or OR4_24(I7979,g6015,g6212,g4950,g4877);
  or OR2_164(g5531,g5349,g3275);
  or OR2_165(g5458,g3466,g5311);
  or OR2_166(g6795,g4867,g6772);
  or OR2_167(g4936,g4827,g4828);
  or OR2_168(g5074,g4792,g4598);
  or OR2_169(g5474,g5363,g5146);
  or OR2_170(g6926,g6798,g6923);
  or OR3_10(g6754,g6676,g6625,g6737);
  or OR2_171(g6273,g5681,g5955);
  or OR2_172(g6444,g6338,g5936);
  or OR4_25(I8378,g5173,g5166,g5235,g5245);
  or OR4_26(I8135,g6194,g5958,g5975,g5997);
  or OR3_11(g5326,g5069,g4410,g3012);
  or OR3_12(I9066,g5189,g5269,g6400);
  or OR2_173(g6927,g6799,g6924);
  or OR2_174(g3751,g3375,g2807);
  or OR2_175(g6660,g6640,g6637);
  or OR2_176(g6679,g6637,g6558);
  or OR4_27(I8208,g6194,g5958,g5975,g5997);
  or OR2_177(g6182,g6047,g6034);
  or OR3_13(g5327,g5077,g4416,g3028);
  or OR2_178(g3743,g3344,g2758);
  or OR2_179(g3856,g3686,g3157);
  or OR2_180(g5303,g5053,g4768);
  or OR2_181(g5696,g5637,g5484);
  or OR2_182(g3992,g1555,g3559);
  or OR2_183(g5472,g5361,g5144);
  or OR2_184(g3863,g3692,g3172);
  or OR2_185(g6437,g6302,g6121);
  or OR2_186(g6917,g6909,g6910);
  or OR2_187(g3857,g3687,g3161);
  or OR2_188(g5533,g5351,g3290);
  or OR2_189(g5697,g5646,g5485);
  or OR2_190(g5013,g4826,g4621);
  or OR2_191(g4627,g4333,g3603);
  or OR2_192(g6454,g6344,g5949);
  or OR2_193(g6296,g6247,g6088);
  or OR2_194(g4646,g4353,g3635);
  or OR4_28(I8138,g4980,g4915,g5025,g5054);
  or OR2_195(g6189,g6060,g6035);
  or OR2_196(g3977,g3653,g3113);
  or OR4_29(I9058,g6156,g6331,g5190,g5164);
  or OR2_197(g6787,g3758,g6766);
  or OR2_198(g5060,g3491,g4819);
  or OR2_199(g6297,g6248,g6089);
  or OR2_200(g3999,g3699,g3181);
  or OR2_201(g6684,g6250,g6643);
  or OR4_30(I7978,g6194,g5958,g5975,g5997);
  or OR2_202(g6109,g5900,g5599);
  or OR2_203(g6791,g6768,g3307);
  or OR2_204(g6309,g6265,g6098);
  or OR2_205(g3732,g3324,g2732);
  or OR2_206(g3533,g3154,g3166);
  or OR4_31(I8385,g6316,g6128,g6131,g6149);
  or OR2_207(g6268,g5677,g5951);
  or OR2_208(g3820,g3287,g2671);
  or OR2_209(g6452,g6342,g5942);
  or OR2_210(g5626,g5496,g3285);
  or OR2_211(g4656,g4369,g3662);
  or OR2_212(g6185,g6055,g5995);
  or OR2_213(g3739,g3334,g2746);
  or OR4_32(I7989,g5202,g4993,g4967,g4980);
  or OR2_214(g3995,g3690,g3170);
  or OR4_33(I8369,g5165,g5159,g5233,g5240);
  or OR4_34(I7971,g5202,g4993,g4967,g4980);
  or OR2_215(g5627,g5497,g3286);
  or OR3_14(g6682,g6478,g6624,g6623);
  or OR2_216(g3942,g3215,g3575);
  or OR2_217(g5583,g5569,g4020);
  or OR2_218(g6173,g6066,g6043);
  or OR2_219(g3954,g3484,g3489);
  or OR2_220(g6920,g6915,g6916);
  or OR2_221(g6261,g5673,g5944);
  or OR2_222(g6793,g6771,g3323);
  or OR2_223(g4948,g4834,g4836);
  or OR2_224(g6246,g5665,g5937);
  or OR2_225(g5224,g5123,g3630);
  or OR2_226(g5277,g5023,g4763);
  or OR2_227(g4438,g4363,g4037);
  or OR2_228(g4773,g4495,g4220);
  or OR2_229(g6689,g6266,g6648);
  or OR2_230(g3998,g3698,g3180);
  or OR4_35(I8774,g6655,g6653,g6651,g6649);
  or OR2_231(g3850,g3680,g3145);
  or OR2_232(g6108,g5898,g5598);
  or OR3_15(g6758,g6673,g6628,g6738);
  or OR2_233(g2896,g2323,g1763);
  or OR2_234(g6455,g6345,g5952);
  or OR2_235(g3986,g3667,g3133);
  or OR2_236(g6846,g5860,g6834);
  or OR2_237(g3503,g3122,g3132);
  or OR4_36(I7969,g6194,g5958,g5975,g5997);
  or OR2_238(g4941,g4829,g4832);
  or OR2_239(g6290,g6245,g6086);
  or OR2_240(g3987,g3669,g3134);
  or OR2_241(g6847,g5861,g6837);
  or OR2_242(g6685,g6256,g6644);
  or OR2_243(g5295,g5047,g4766);
  or OR2_244(g4473,g3575,g4253);
  or OR2_245(g3991,g3685,g3156);
  or OR4_37(I7988,g6015,g6212,g4950,g4877);
  or OR2_246(g5471,g5360,g5143);
  or OR4_38(I8368,g6148,g6321,g5176,g5184);
  or OR2_247(g6257,g5671,g5941);
  or OR2_248(g6301,g6254,g6092);
  or OR4_39(g6673,g6559,g6640,g4416,g2950);
  or OR4_40(I8080,g6015,g6212,g4950,g4877);
  or OR2_249(g6669,g6613,g4679);
  or OR2_250(g3877,g3651,g3659);
  or OR4_41(I8126,g6194,g5958,g5975,g5997);
  or OR2_251(g5062,g4661,g4666);
  or OR2_252(g6480,I8360,g6359);
  or OR4_42(I8779,g6605,g6656,g6654,g6652);
  or OR2_253(g6688,g6263,g6647);
  or OR2_254(g5085,g4694,g4280);
  or OR2_255(I7981,g4915,g5025);
  or OR4_43(I8127,g6015,g6212,g4950,g4877);
  or OR2_256(g4433,g4354,g4032);
  or OR4_44(I8346,g6159,g6334,g5163,g5191);
  or OR2_257(g5812,g5376,g5618);
  or OR2_258(g4859,g4730,g4486);
  or OR2_259(g6665,I8778,I8779);
  or OR2_260(g5473,g5362,g5145);
  or OR4_45(I8347,g5188,g5157,g5154,g5193);
  or OR2_261(g6303,g6258,g6094);
  or OR2_262(g5069,g1595,g4688);
  or OR4_46(I9064,g6323,g6829,g6831,g6155);
  or OR2_263(g4497,g4166,g3784);
  or OR4_47(I8210,g5202,g4993,g4967,g4980);
  or OR2_264(g5377,g5217,g4949);
  or OR2_265(g3837,g3609,g3613);
  or OR2_266(g6116,g5910,g5617);
  or OR4_48(I8117,g6194,g5958,g5975,g5997);
  or OR2_267(g4001,g3702,g3190);
  or OR2_268(g3842,g3670,g3135);
  or OR2_269(g5291,g5043,g4764);
  or OR2_270(g3941,g3479,g2873);
  or OR2_271(g5694,g5633,g5482);
  or OR2_272(g6936,g5438,g6935);
  or OR2_273(g4068,g3293,g2685);
  or OR4_49(I8079,g6194,g5958,g5975,g5997);
  or OR2_274(g4468,g4214,g3831);
  or OR2_275(g4866,g4756,g4491);
  or OR2_276(g3829,g3294,g3305);
  or OR4_50(I8356,g6311,g6123,g6125,g6141);
  or OR2_277(g3733,g3325,g2733);
  or OR2_278(g6937,g4616,g6934);
  or OR2_279(g6479,I8349,g6335);
  or OR2_280(g6294,g6249,g6090);
  or OR2_281(g5065,g4667,g4671);
  or OR2_282(g5228,g5096,g4800);
  or OR4_51(I8357,g6145,g6318,g5171,g5187);
  or OR2_283(g3849,g3618,g3625);
  or OR2_284(g6704,g6660,g492);
  or OR2_285(g4599,g3499,g4230);
  or OR2_286(g6453,g6343,g5945);
  or OR2_287(g4544,g4410,g2995);
  or OR4_52(I8778,g6612,g6611,g6609,g6607);
  or OR2_288(g2924,g2095,g1573);
  or OR2_289(g4427,g4373,g3668);
  or OR2_290(g4446,g4383,g4043);
  or OR2_291(g3870,g3700,g3182);
  or OR3_16(g6683,g6465,g6622,g6621);
  or OR2_292(g5676,g5559,g5424);
  or OR2_293(g4637,g4344,g3619);
  or OR2_294(g3972,g3646,g3103);
  or OR2_295(g6782,g6719,g6749);
  or OR2_296(g6661,I8773,I8774);
  or OR2_297(g4757,g4456,g4158);
  or OR2_298(g6292,g6243,g6084);
  or OR2_299(g4811,g4429,g4432);
  or OR2_300(g4642,g4348,g3628);
  or OR2_301(g4447,g4384,g4044);
  or OR2_302(g5624,g5494,g3280);
  or OR2_303(g5068,g4673,g4677);
  or OR2_304(g4654,g4362,g3654);
  or OR2_305(g3891,g3683,g3688);
  or OR2_306(g3913,g3449,g2860);
  or OR2_307(I7990,g4915,g5025);
  or OR2_308(g6702,g6659,g496);
  or OR2_309(g6919,g6912,g6914);
  or OR2_310(I8120,g4915,g5025);
  or OR2_311(g4243,g4053,g4058);
  or OR2_312(g5699,g5660,g5487);
  or OR2_313(g5241,g5069,g2067);
  or OR2_314(g4234,g3921,g478);
  or OR2_315(g3815,g3282,g2659);
  or OR2_316(g5386,g5227,g669);
  or OR2_317(g6789,g3764,g6769);
  or OR4_53(I8082,g4980,g4915,g5025,g5054);
  or OR2_318(g5370,g5211,g4937);
  or OR2_319(g3828,g3304,g1351);
  or OR4_54(I9065,g6158,g6333,g5152,g5156);
  or OR2_320(g3746,g3357,g2771);
  or OR2_321(g5083,g4688,g4271);
  or OR2_322(g6907,g6874,g3358);
  or OR2_323(g5622,g5492,g3277);
  or OR2_324(g6690,g6270,g6650);
  or OR4_55(g6482,I8376,I8377,I8378,I8379);
  or OR2_325(g4652,g4358,g3645);
  or OR2_326(g4549,g4416,g3013);
  or OR2_327(g3747,g3365,g2781);
  or OR2_328(g3855,g3626,g3631);
  or OR2_329(g5695,g5635,g5483);
  or OR2_330(g6110,g5883,g5996);
  or OR2_331(g6310,g6269,g6099);
  or OR2_332(g5016,g4789,g4592);
  or OR3_17(g6762,g6679,g6628,g6739);
  or OR2_333(g4740,g4448,g4154);
  or OR4_56(I8394,g6154,g6329,g5186,g5172);
  or OR2_334(g6556,g6339,g6467);
  or OR2_335(g6930,g6740,g6928);
  or OR2_336(g3599,g2935,g1637);
  or OR2_337(g3821,g2951,g3466);
  or OR2_338(g4860,g4735,g4488);
  or OR2_339(g6237,g5912,g2381);
  or OR2_340(g4645,g4352,g3633);
  or OR3_18(g6844,I9057,I9058,I9059);
  or OR4_57(I8773,g6610,g6608,g6606,g6604);
  or OR2_341(g5629,g5499,g3298);
  or OR2_342(g4607,g4232,g3899);
  or OR2_343(g6705,g6693,g4835);
  or OR2_344(g5800,g5369,g5600);
  or OR2_345(g6242,g2356,g6075);
  or OR2_346(g3841,g3614,g3617);
  or OR2_347(g6918,g6911,g6913);
  or OR2_348(g5348,g5317,g5122);
  or OR2_349(g3858,g3629,g3636);
  or OR2_350(g5698,g5648,g5486);
  or OR2_351(g4630,g4339,g3610);
  or OR2_352(g6921,g6908,g6816);
  or OR2_353(g5367,g5199,g4928);
  nand NAND3_0(g1777,g1060,g102,g89);
  nand NAND2_0(I7217,g152,I7216);
  nand NAND2_1(I7571,g5678,I7569);
  nand NAND4_0(g5686,g5546,g1017,g1551,g2916);
  nand NAND2_2(I2073,g15,I2072);
  nand NAND2_3(I2796,g804,I2795);
  nand NAND2_4(g948,I2014,I2015);
  nand NAND2_5(I4205,g743,I4203);
  nand NAND2_6(I3875,g285,I3874);
  nand NAND3_1(g3330,g1815,g1797,g3109);
  nand NAND2_7(g4151,I5536,I5537);
  nand NAND3_2(g2435,g1138,g1777,g1157);
  nand NAND2_8(I5658,g3983,I5657);
  nand NAND2_9(g1558,I2527,I2528);
  nand NAND2_10(I4444,g2092,g606);
  nand NAND2_11(I5271,g3710,I5269);
  nand NAND2_12(I2898,g1027,I2897);
  nand NAND2_13(I2797,g798,I2795);
  nand NAND2_14(I2245,g567,I2244);
  nand NAND2_15(I3988,g291,g2544);
  nand NAND2_16(g1574,I2543,I2544);
  nand NAND4_1(g3529,g3200,g2215,g2976,g2968);
  nand NAND2_17(I1963,g242,I1961);
  nand NAND2_18(I5209,g3271,I5207);
  nand NAND2_19(I7562,g74,g5676);
  nand NAND2_20(g5506,I7231,I7232);
  nand NAND2_21(g5111,I6744,I6745);
  nand NAND2_22(I4182,g2292,g749);
  nand NAND2_23(I6186,g4301,I6185);
  nand NAND2_24(I7441,g594,I7439);
  nand NAND2_25(I6026,g4223,g4221);
  nand NAND2_26(I2768,g743,I2766);
  nand NAND2_27(I3933,g288,g2473);
  nand NAND3_3(g5853,g5638,g2053,g1076);
  nand NAND2_28(g2731,I3894,I3895);
  nand NAND2_29(g5507,I7238,I7239);
  nand NAND2_30(g2966,I4160,I4161);
  nand NAND2_31(I2934,g1436,I2933);
  nand NAND2_32(I3179,g736,I3177);
  nand NAND2_33(I6187,g3955,I6185);
  nand NAND2_34(I6027,g4223,I6026);
  nand NAND3_4(g2009,g901,g1387,g905);
  nand NAND2_35(I4233,g2267,g798);
  nand NAND2_36(g2769,I3953,I3954);
  nand NAND2_37(g1044,I2081,I2082);
  nand NAND4_2(g4674,g4550,g1514,g2107,g2897);
  nand NAND2_38(I7569,g79,g5678);
  nand NAND2_39(I6391,g4504,I6390);
  nand NAND4_3(g3525,g3192,g3002,g2197,g2179);
  nand NAND4_4(g4680,g4550,g1514,g1006,g2897);
  nand NAND2_40(I2081,g25,I2080);
  nand NAND2_41(I8195,g471,I8194);
  nand NAND2_42(g1534,I2498,I2499);
  nand NAND2_43(I2497,g1042,g1036);
  nand NAND2_44(g939,I1987,I1988);
  nand NAND2_45(I5269,g3705,g3710);
  nand NAND3_5(g3985,g1138,g3718,g2142);
  nand NAND2_46(g1036,I2061,I2062);
  nand NAND2_47(I2676,g131,I2674);
  nand NAND2_48(g1749,I2767,I2768);
  nand NAND2_49(g6097,g2954,g5857);
  nand NAND3_6(g6783,g6747,g5068,g5066);
  nand NAND2_50(g5776,I7528,I7529);
  nand NAND2_51(I7434,g5554,I7432);
  nand NAND2_52(g1042,I2073,I2074);
  nand NAND2_53(I7210,g5367,I7208);
  nand NAND4_5(g3530,g3204,g3023,g2197,g2179);
  nand NAND2_54(I6964,g586,I6962);
  nand NAND2_55(I5208,g3267,I5207);
  nand NAND2_56(I5302,g3505,I5300);
  nand NAND2_57(g5777,I7535,I7536);
  nand NAND2_58(g4613,I6195,I6196);
  nand NAND2_59(I2544,g774,I2542);
  nand NAND2_60(g1138,g102,g98);
  nand NAND2_61(I1994,g504,g218);
  nand NAND2_62(I4445,g2092,I4444);
  nand NAND2_63(I2061,g7,I2060);
  nand NAND2_64(I5189,g3593,I5187);
  nand NAND2_65(g4903,g4717,g858);
  nand NAND2_66(I3178,g1706,I3177);
  nand NAND2_67(I4920,g3522,I4919);
  nand NAND2_68(g2951,g2142,g1797);
  nand NAND4_6(g3518,g3177,g3023,g3007,g2981);
  nand NAND2_69(I2003,g500,g212);
  nand NAND3_7(g6717,g6669,g5065,g5062);
  nand NAND2_70(I3916,g2449,I3914);
  nand NAND4_7(g5864,g5649,g1529,g1088,g2068);
  nand NAND3_8(g2008,g866,g873,g1784);
  nand NAND2_71(I5309,g3512,I5307);
  nand NAND2_72(I7432,g111,g5554);
  nand NAND2_73(I4203,g2255,g743);
  nand NAND4_8(g3521,g3187,g3023,g3007,g2179);
  nand NAND2_74(I5759,g3836,g3503);
  nand NAND2_75(I6962,g4874,g586);
  nand NAND2_76(I6659,g4762,g3541);
  nand NAND2_77(I4940,g3437,I4939);
  nand NAND2_78(I2935,g345,I2933);
  nand NAND2_79(g2266,I3412,I3413);
  nand NAND2_80(I2542,g821,g774);
  nand NAND2_81(I3412,g1419,I3411);
  nand NAND2_82(I3189,g1716,I3188);
  nand NAND2_83(g5634,g5563,g4767);
  nand NAND2_84(I3990,g2544,I3988);
  nand NAND2_85(g2960,I4151,I4152);
  nand NAND2_86(g5926,g5741,g639);
  nand NAND4_9(g3511,g3158,g3002,g2976,g2968);
  nand NAND2_87(I7439,g5515,g594);
  nand NAND2_88(I2090,g33,I2089);
  nand NAND4_10(g5862,g5649,g1529,g1535,g2068);
  nand NAND2_89(I9050,g6832,g3598);
  nand NAND2_90(I5766,g3961,g3957);
  nand NAND3_9(g1582,g784,g774,g821);
  nand NAND2_91(g1793,g94,g1084);
  nand NAND2_92(g3968,I5227,I5228);
  nand NAND2_93(I7527,g49,g5662);
  nand NAND2_94(I5226,g3259,g3263);
  nand NAND2_95(g4049,g3677,g3425);
  nand NAND2_96(I7224,g161,I7223);
  nand NAND2_97(I5767,g3961,I5766);
  nand NAND2_98(I5535,g3907,g654);
  nand NAND2_99(I5227,g3259,I5226);
  nand NAND2_100(g5947,g5821,g2944);
  nand NAND2_101(g3742,I4920,I4921);
  nand NAND4_11(g5873,g5649,g1017,g1564,g2113);
  nand NAND2_102(g4504,I6027,I6028);
  nand NAND2_103(I7244,g188,g5377);
  nand NAND3_10(g5869,g5649,g1076,g2081);
  nand NAND2_104(I5188,g3589,I5187);
  nand NAND2_105(g3983,I5270,I5271);
  nand NAND4_12(g4678,g2897,g2101,g1514,g4550);
  nand NAND2_106(g6843,I9051,I9052);
  nand NAND2_107(g3961,I5208,I5209);
  nand NAND2_108(I5308,g478,I5307);
  nand NAND2_109(I2506,g1047,g1044);
  nand NAND2_110(I3445,g1689,g729);
  nand NAND2_111(g2061,I3169,I3170);
  nand NAND2_112(I3169,g1540,I3168);
  nand NAND3_11(g6740,g6703,g6457,g4936);
  nand NAND2_113(I7556,g69,I7555);
  nand NAND2_114(g4007,I5308,I5309);
  nand NAND2_115(I5196,g3567,I5195);
  nand NAND2_116(I7563,g74,I7562);
  nand NAND2_117(g5684,I7440,I7441);
  nand NAND2_118(I2507,g1047,I2506);
  nand NAND2_119(I1995,g504,I1994);
  nand NAND2_120(g2307,I3446,I3447);
  nand NAND2_121(I7237,g179,g5374);
  nand NAND2_122(g2858,g1815,g2577);
  nand NAND2_123(g2757,I3934,I3935);
  nand NAND2_124(I6744,g4708,I6743);
  nand NAND2_125(I4183,g2292,I4182);
  nand NAND2_126(I7557,g5674,I7555);
  nand NAND2_127(I2300,g830,I2299);
  nand NAND2_128(I3188,g1716,g791);
  nand NAND4_13(g5865,g5649,g1088,g1076,g2068);
  nand NAND2_129(I5197,g3571,I5195);
  nand NAND2_130(I4161,g619,I4159);
  nand NAND2_131(I3741,g349,I3739);
  nand NAND2_132(g5019,I6660,I6661);
  nand NAND2_133(I5257,g3714,g3719);
  nand NAND4_14(g3532,g3212,g2215,g3007,g2981);
  nand NAND2_134(I2528,g719,I2526);
  nand NAND2_135(I5301,g471,I5300);
  nand NAND2_136(g1743,g1064,g94);
  nand NAND2_137(g1411,g314,g873);
  nand NAND2_138(g3012,I4204,I4205);
  nand NAND2_139(g5504,I7217,I7218);
  nand NAND2_140(I6175,g4236,g571);
  nand NAND2_141(I3455,g1691,g784);
  nand NAND2_142(I6500,g4504,I6499);
  nand NAND3_12(g1573,g729,g719,g766);
  nand NAND2_143(I3846,g284,g2370);
  nand NAND2_144(I4210,g2294,g804);
  nand NAND2_145(g4803,I6474,I6475);
  nand NAND2_146(g3109,g2360,g1064);
  nand NAND2_147(g2698,I3847,I3848);
  nand NAND2_148(g3957,I5196,I5197);
  nand NAND2_149(I6499,g4504,g3541);
  nand NAND4_15(g4816,g996,g4550,g1518,g2073);
  nand NAND2_150(I3847,g284,I3846);
  nand NAND2_151(I7520,g361,g5659);
  nand NAND2_152(I4784,g622,I4782);
  nand NAND2_153(I1952,g524,I1951);
  nand NAND4_16(g3539,g2591,g2215,g2197,g2981);
  nand NAND2_154(I8202,g478,I8201);
  nand NAND2_155(I1986,g508,g224);
  nand NAND2_156(I2933,g1436,g345);
  nand NAND2_157(I5760,g3836,I5759);
  nand NAND2_158(g4301,I5767,I5768);
  nand NAND2_159(I1970,g516,I1969);
  nand NAND2_160(I7225,g5370,I7223);
  nand NAND2_161(I6660,g4762,I6659);
  nand NAND2_162(g5502,I7209,I7210);
  nand NAND2_163(I3168,g1540,g1534);
  nand NAND2_164(I1987,g508,I1986);
  nand NAND2_165(g1316,I2300,I2301);
  nand NAND2_166(I2674,g710,g131);
  nand NAND4_17(g4669,g4550,g1017,g1680,g2897);
  nand NAND2_167(I3411,g1419,g616);
  nand NAND2_168(I7245,g188,I7244);
  nand NAND2_169(g2607,I3740,I3741);
  nand NAND2_170(g5308,I6963,I6964);
  nand NAND2_171(g2311,I3456,I3457);
  nand NAND4_18(g3535,g3216,g2215,g2197,g2968);
  nand NAND2_172(g5455,g2330,g5311);
  nand NAND2_173(I4782,g2846,g622);
  nand NAND2_174(I9052,g3598,I9050);
  nand NAND2_175(I3126,g1279,I3125);
  nand NAND2_176(I3400,g135,I3398);
  nand NAND2_177(I4526,g2909,g646);
  nand NAND2_178(g5780,I7556,I7557);
  nand NAND2_179(g3246,I4527,I4528);
  nand NAND3_13(g3502,g1411,g1402,g2795);
  nand NAND2_180(g4608,I6176,I6177);
  nand NAND2_181(I4919,g3522,g650);
  nand NAND3_14(g2100,g1588,g804,g791);
  nand NAND2_182(I7230,g170,g5372);
  nand NAND2_183(I7433,g111,I7432);
  nand NAND2_184(I3127,g1276,I3125);
  nand NAND2_185(g3028,I4234,I4235);
  nand NAND2_186(I2795,g804,g798);
  nand NAND2_187(I5784,g628,I5782);
  nand NAND2_188(I4527,g2909,I4526);
  nand NAND2_189(I7550,g5672,I7548);
  nand NAND2_190(I4546,g2853,I4545);
  nand NAND2_191(I6745,g582,I6743);
  nand NAND2_192(I5294,g625,I5292);
  nand NAND2_193(I6963,g4874,I6962);
  nand NAND3_15(g3741,g901,g3433,g2340);
  nand NAND2_194(g1157,g89,g107);
  nand NAND2_195(I2499,g1036,I2497);
  nand NAND2_196(g937,I1979,I1980);
  nand NAND2_197(g4472,g3380,g4253);
  nand NAND3_16(g2010,g1473,g1470,g1459);
  nand NAND2_198(g928,I1962,I1963);
  nand NAND2_199(I7097,g5194,g574);
  nand NAND2_200(I4547,g353,I4545);
  nand NAND2_201(I3697,g1570,g642);
  nand NAND2_202(I3914,g287,g2449);
  nand NAND2_203(I2543,g821,I2542);
  nand NAND2_204(I3413,g616,I3411);
  nand NAND2_205(I7218,g5368,I7216);
  nand NAND2_206(I7312,g5364,I7311);
  nand NAND4_19(g3538,g2588,g2215,g2197,g2179);
  nand NAND2_207(g5505,I7224,I7225);
  nand NAND2_208(g1075,I2109,I2110);
  nand NAND2_209(I2014,g532,I2013);
  nand NAND2_210(g2804,I4009,I4010);
  nand NAND3_17(g6742,g6683,g932,g6716);
  nand NAND2_211(I6185,g4301,g3955);
  nand NAND4_20(g5863,g5649,g1076,g1535,g2068);
  nand NAND2_212(I3739,g2021,g349);
  nand NAND2_213(I2022,g528,I2021);
  nand NAND2_214(I5782,g3810,g628);
  nand NAND2_215(I7576,g84,g5680);
  nand NAND4_21(g5688,g5546,g1585,g2084,g2916);
  nand NAND4_22(g5857,g5638,g1552,g1017,g2062);
  nand NAND2_216(I3190,g791,I3188);
  nand NAND2_217(I5292,g3421,g625);
  nand NAND2_218(g1764,I2796,I2797);
  nand NAND2_219(I3954,g2497,I3952);
  nand NAND2_220(g5779,I7549,I7550);
  nand NAND2_221(I7577,g84,I7576);
  nand NAND2_222(I5647,g3974,g3968);
  nand NAND4_23(g3531,g3209,g2215,g2976,g2179);
  nand NAND2_223(I1980,g230,I1978);
  nand NAND2_224(g5508,I7245,I7246);
  nand NAND2_225(I4150,g2551,g139);
  nand NAND2_226(g6873,g6848,g3621);
  nand NAND2_227(g6095,g2952,g5854);
  nand NAND2_228(I4009,g292,I4008);
  nand NAND2_229(I2675,g710,I2674);
  nand NAND2_230(g926,I1952,I1953);
  nand NAND2_231(I3894,g286,I3893);
  nand NAND2_232(I4212,g804,I4210);
  nand NAND2_233(g5565,I7312,I7313);
  nand NAND2_234(I6028,g4221,I6026);
  nand NAND2_235(I2109,g602,I2108);
  nand NAND2_236(I5244,g3247,I5242);
  nand NAND3_18(g1402,g310,g866,g873);
  nand NAND2_237(I4921,g650,I4919);
  nand NAND2_238(I7536,g5666,I7534);
  nand NAND2_239(I7223,g161,g5370);
  nand NAND2_240(I2498,g1042,I2497);
  nand NAND2_241(I1951,g524,g248);
  nand NAND2_242(I7522,g5659,I7520);
  nand NAND2_243(I3952,g289,g2497);
  nand NAND2_244(g5775,I7521,I7522);
  nand NAND2_245(I8201,g478,g6192);
  nand NAND2_246(g2024,I3126,I3127);
  nand NAND2_247(g2795,g1997,g866);
  nand NAND2_248(g4004,I5301,I5302);
  nand NAND2_249(I6196,g631,I6194);
  nand NAND2_250(I3970,g290,g2518);
  nand NAND2_251(I4941,g357,I4939);
  nand NAND2_252(I5657,g3983,g3979);
  nand NAND2_253(I7542,g59,I7541);
  nand NAND2_254(I2897,g1027,g634);
  nand NAND2_255(I2682,g918,I2681);
  nand NAND2_256(I2766,g749,g743);
  nand NAND2_257(g3013,I4211,I4212);
  nand NAND2_258(I5242,g3242,g3247);
  nand NAND2_259(I7529,g5662,I7527);
  nand NAND2_260(g1822,g1070,g1084);
  nand NAND2_261(I3876,g2397,I3874);
  nand NAND2_262(I2091,g29,I2089);
  nand NAND2_263(I3915,g287,I3914);
  nand NAND2_264(I9051,g6832,I9050);
  nand NAND2_265(I2767,g749,I2766);
  nand NAND2_266(I1979,g512,I1978);
  nand NAND2_267(g3597,I4783,I4784);
  nand NAND3_19(g2831,g2007,g862,g1784);
  nand NAND2_268(g5683,I7433,I7434);
  nand NAND2_269(g5778,I7542,I7543);
  nand NAND2_270(I2015,g260,I2013);
  nand NAND2_271(g930,I1970,I1971);
  nand NAND2_272(g5782,I7570,I7571);
  nand NAND2_273(g4002,I5293,I5294);
  nand NAND2_274(I2246,g598,I2244);
  nand NAND2_275(I6743,g4708,g582);
  nand NAND2_276(I7549,g64,I7548);
  nand NAND2_277(g2947,g1411,g2026);
  nand NAND2_278(g4762,I6391,I6392);
  nand NAND3_20(g2095,g1584,g749,g736);
  nand NAND2_279(g944,I2004,I2005);
  nand NAND2_280(I6474,g4541,I6473);
  nand NAND2_281(I7232,g5372,I7230);
  nand NAND2_282(I1953,g248,I1951);
  nand NAND2_283(g2719,I3875,I3876);
  nand NAND2_284(I8203,g6192,I8201);
  nand NAND2_285(I4008,g292,g2568);
  nand NAND2_286(g4237,g4049,g4017);
  nand NAND2_287(g1829,I2898,I2899);
  nand NAND2_288(g901,g314,g310);
  nand NAND2_289(g941,I1995,I1996);
  nand NAND2_290(I7570,g79,I7569);
  nand NAND2_291(I2108,g602,g610);
  nand NAND2_292(g1540,I2507,I2508);
  nand NAND4_24(g4814,g4550,g1575,g1550,g2073);
  nand NAND2_293(I7311,g5364,g590);
  nand NAND2_294(I5270,g3705,I5269);
  nand NAND2_295(g2745,I3915,I3916);
  nand NAND3_21(g1797,g98,g1064,g1070);
  nand NAND2_296(g2791,I3989,I3990);
  nand NAND2_297(I7239,g5374,I7237);
  nand NAND4_25(g3526,g3196,g3023,g2197,g2981);
  nand NAND3_22(g6741,g6705,g6461,g4941);
  nand NAND2_298(I8196,g6188,I8194);
  nand NAND2_299(I3895,g2422,I3893);
  nand NAND2_300(I4783,g2846,I4782);
  nand NAND2_301(I2021,g528,g254);
  nand NAND2_302(g905,g301,g319);
  nand NAND2_303(g3276,I4546,I4547);
  nand NAND2_304(g6774,g6754,g6750);
  nand NAND2_305(I5207,g3267,g3271);
  nand NAND2_306(I2301,g341,I2299);
  nand NAND2_307(I5259,g3719,I5257);
  nand NAND2_308(I7440,g5515,I7439);
  nand NAND2_309(I7528,g49,I7527);
  nand NAND2_310(g4640,g4402,g1056);
  nand NAND4_26(g4812,g4550,g1560,g1559,g2073);
  nand NAND2_311(g1845,I2934,I2935);
  nand NAND2_312(g6397,I8202,I8203);
  nand NAND2_313(I5768,g3957,I5766);
  nand NAND2_314(I1978,g512,g230);
  nand NAND2_315(g4610,I6186,I6187);
  nand NAND2_316(I5228,g3263,I5226);
  nand NAND2_317(I2074,g11,I2072);
  nand NAND3_23(g3140,g2409,g1060,g1620);
  nand NAND2_318(I6390,g4504,g4610);
  nand NAND2_319(I3177,g1706,g736);
  nand NAND2_320(I4152,g139,I4150);
  nand NAND2_321(I6501,g3541,I6499);
  nand NAND2_322(I7548,g64,g5672);
  nand NAND2_323(g1815,g102,g1070);
  nand NAND2_324(I7555,g69,g5674);
  nand NAND4_27(g3517,g3173,g3002,g2976,g2179);
  nand NAND2_325(I2080,g25,g19);
  nand NAND2_326(I4211,g2294,I4210);
  nand NAND2_327(I3399,g1826,I3398);
  nand NAND2_328(I5195,g3567,g3571);
  nand NAND2_329(I7313,g590,I7311);
  nand NAND2_330(g2582,I3698,I3699);
  nand NAND2_331(I4939,g3437,g357);
  nand NAND2_332(g950,I2022,I2023);
  nand NAND2_333(g4819,I6500,I6501);
  nand NAND2_334(I7521,g361,I7520);
  nand NAND2_335(I2023,g254,I2021);
  nand NAND2_336(I4446,g606,I4444);
  nand NAND2_337(I5783,g3810,I5782);
  nand NAND2_338(g2940,g197,g2381);
  nand NAND2_339(g4825,g4472,g4465);
  nand NAND2_340(I5293,g3421,I5292);
  nand NAND2_341(I5761,g3503,I5759);
  nand NAND2_342(I1971,g236,I1969);
  nand NAND2_343(I3972,g2518,I3970);
  nand NAND2_344(I4159,g2015,g619);
  nand NAND2_345(I6661,g3541,I6659);
  nand NAND2_346(g1398,g306,g889);
  nand NAND2_347(I6475,g578,I6473);
  nand NAND2_348(I3934,g288,I3933);
  nand NAND2_349(I7541,g59,g5669);
  nand NAND2_350(I2508,g1044,I2506);
  nand NAND4_28(g5854,g5638,g1683,g1552,g2062);
  nand NAND2_351(g4465,g319,g4253);
  nand NAND2_352(I2072,g15,g11);
  nand NAND2_353(I7238,g179,I7237);
  nand NAND2_354(g3955,I5188,I5189);
  nand NAND2_355(I7209,g143,I7208);
  nand NAND2_356(g5431,I7098,I7099);
  nand NAND2_357(I2681,g918,g613);
  nand NAND2_358(I2013,g532,g260);
  nand NAND2_359(I4234,g2267,I4233);
  nand NAND2_360(g2780,I3971,I3972);
  nand NAND2_361(g2067,I3178,I3179);
  nand NAND2_362(I1962,g520,I1961);
  nand NAND2_363(I5258,g3714,I5257);
  nand NAND3_24(g1387,g862,g314,g301);
  nand NAND2_364(I2060,g7,g3);
  nand NAND2_365(g5781,I7563,I7564);
  nand NAND2_366(g2263,I3399,I3400);
  nand NAND2_367(g4221,I5648,I5649);
  nand NAND2_368(g1359,g866,g306);
  nand NAND2_369(I7231,g170,I7230);
  nand NAND2_370(I3953,g289,I3952);
  nand NAND2_371(I5187,g3589,g3593);
  nand NAND3_25(g5852,g5638,g2053,g1661);
  nand NAND4_29(g3520,g3183,g3002,g2197,g2968);
  nand NAND2_372(g1047,I2090,I2091);
  nand NAND2_373(I7099,g574,I7097);
  nand NAND2_374(I3848,g2370,I3846);
  nand NAND2_375(I3699,g642,I3697);
  nand NAND2_376(I3398,g1826,g135);
  nand NAND2_377(I1969,g516,g236);
  nand NAND2_378(I5307,g478,g3512);
  nand NAND2_379(g3974,I5243,I5244);
  nand NAND2_380(I5536,g3907,I5535);
  nand NAND2_381(g1417,g873,g889);
  nand NAND2_382(I7543,g5669,I7541);
  nand NAND2_383(g5943,g5818,g2940);
  nand NAND2_384(I7534,g54,g5666);
  nand NAND2_385(g4319,I5783,I5784);
  nand NAND2_386(I3893,g286,g2422);
  nand NAND2_387(g2080,I3189,I3190);
  nand NAND2_388(I2683,g613,I2681);
  nand NAND2_389(I5537,g654,I5535);
  nand NAND2_390(I3170,g1534,I3168);
  nand NAND2_391(I3125,g1279,g1276);
  nand NAND2_392(I5243,g3242,I5242);
  nand NAND2_393(I1988,g224,I1986);
  nand NAND2_394(I6194,g4199,g631);
  nand NAND2_395(g3207,I4445,I4446);
  nand NAND2_396(I2526,g766,g719);
  nand NAND2_397(g6929,g4536,g6927);
  nand NAND2_398(g3215,g2340,g1402);
  nand NAND2_399(I3446,g1689,I3445);
  nand NAND2_400(I7208,g143,g5367);
  nand NAND2_401(g5783,I7577,I7578);
  nand NAND2_402(I4545,g2853,g353);
  nand NAND2_403(I2004,g500,I2003);
  nand NAND2_404(I2527,g766,I2526);
  nand NAND2_405(I5649,g3968,I5647);
  nand NAND2_406(g6778,g6762,g6758);
  nand NAND2_407(g1686,I2675,I2676);
  nand NAND2_408(g4223,I5658,I5659);
  nand NAND2_409(I1996,g218,I1994);
  nand NAND2_410(I3447,g729,I3445);
  nand NAND2_411(I4204,g2255,I4203);
  nand NAND2_412(I3874,g285,g2397);
  nand NAND2_413(g2944,g269,g2381);
  nand NAND2_414(g1253,I2245,I2246);
  nand NAND3_26(g2434,g1064,g1070,g1620);
  nand NAND2_415(I2299,g830,g341);
  nand NAND3_27(g5866,g5649,g1529,g2081);
  nand NAND2_416(g1687,I2682,I2683);
  nand NAND2_417(I3935,g2473,I3933);
  nand NAND2_418(g4017,g107,g3425);
  nand NAND2_419(I4528,g646,I4526);
  nand NAND2_420(I2244,g567,g598);
  nand NAND2_421(I4151,g2551,I4150);
  nand NAND2_422(I6392,g4610,I6390);
  nand NAND2_423(I4010,g2568,I4008);
  nand NAND2_424(I2082,g19,I2080);
  nand NAND4_30(g5818,g5638,g2056,g1666,g1661);
  nand NAND2_425(g3979,I5258,I5259);
  nand NAND2_426(I6176,g4236,I6175);
  nand NAND2_427(I4235,g798,I4233);
  nand NAND2_428(I2110,g610,I2108);
  nand NAND2_429(I7098,g5194,I7097);
  nand NAND2_430(I3456,g1691,I3455);
  nand NAND4_31(g5821,g5638,g2056,g1076,g1666);
  nand NAND2_431(I3698,g1570,I3697);
  nand NAND2_432(g2995,I4183,I4184);
  nand NAND2_433(I6473,g4541,g578);
  nand NAND2_434(I5659,g3979,I5657);
  nand NAND2_435(g5636,g5564,g4769);
  nand NAND2_436(I6177,g571,I6175);
  nand NAND2_437(I2899,g634,I2897);
  nand NAND2_438(I3457,g784,I3455);
  nand NAND2_439(I3989,g291,I3988);
  nand NAND2_440(I3971,g290,I3970);
  nand NAND2_441(I4160,g2015,I4159);
  nand NAND2_442(I2089,g33,g29);
  nand NAND2_443(g4670,g4611,g3528);
  nand NAND4_32(g4813,g4550,g965,g1560,g2073);
  nand NAND2_444(I3740,g2021,I3739);
  nand NAND2_445(I8194,g471,g6188);
  nand NAND2_446(I5300,g471,g3505);
  nand NAND3_28(g3893,g3664,g3656,g3647);
  nand NAND2_447(g6928,g4532,g6926);
  nand NAND2_448(I7578,g5680,I7576);
  nand NAND2_449(I7535,g54,I7534);
  nand NAND2_450(I1961,g520,g242);
  nand NAND4_33(g3544,g2594,g2215,g2197,g2179);
  nand NAND2_451(g6394,I8195,I8196);
  nand NAND2_452(I5648,g3974,I5647);
  nand NAND2_453(I7246,g5377,I7244);
  nand NAND2_454(g3756,I4940,I4941);
  nand NAND2_455(I2062,g3,I2060);
  nand NAND2_456(I6195,g4199,I6194);
  nand NAND2_457(I7216,g152,g5368);
  nand NAND4_34(g3536,g3219,g2215,g3007,g2179);
  nand NAND2_458(I7564,g5676,I7562);
  nand NAND2_459(g4300,I5760,I5761);
  nand NAND2_460(I4184,g749,I4182);
  nand NAND2_461(I2005,g212,I2003);
  nand NAND2_462(g5318,g676,g5060);
  nand NAND4_35(g5872,g5649,g1557,g1564,g2113);
  nor NOR2_0(g5552,g5354,g5356);
  nor NOR2_1(g4235,g3780,g3362);
  nor NOR2_2(g6073,g197,g5862);
  nor NOR2_3(g4776,g4449,g4453);
  nor NOR2_4(g4777,g4457,g4459);
  nor NOR2_5(g4238,g3755,g3279);
  nor NOR4_0(g6433,g6385,g3733,g4092,g4314);
  nor NOR2_6(g6496,g952,g6354);
  nor NOR2_7(g1422,g1039,g913);
  nor NOR2_8(g3931,g3353,g3361);
  nor NOR2_9(g1560,g996,g980);
  nor NOR2_10(g3905,g3512,g478);
  nor NOR2_11(g5094,g4685,g4686);
  nor NOR2_12(g3973,g3368,g3374);
  nor NOR2_13(g3528,g1802,g3167);
  nor NOR2_14(g5541,g5388,g1880);
  nor NOR2_15(g3621,g1407,g2842);
  nor NOR2_16(g1449,g489,g1048);
  nor NOR2_17(g3965,g3359,g3367);
  nor NOR2_18(g3933,g3327,g3336);
  nor NOR4_1(g6280,I7978,I7979,I7980,I7981);
  nor NOR2_19(g2433,g1418,g1449);
  nor NOR3_0(g1470,g937,g930,g928);
  nor NOR4_2(g6427,g6376,g4086,g4074,g4068);
  nor NOR4_3(g6446,g6385,g4334,g4092,g4314);
  nor NOR4_4(g6359,I8135,I8136,I8137,I8138);
  nor NOR3_1(g1459,g926,g950,g948);
  nor NOR2_20(g4584,g4164,g4168);
  nor NOR2_21(g3926,g3338,g3350);
  nor NOR4_5(g6279,I7969,I7970,I7971,I7972);
  nor NOR2_22(g5265,g4863,g4865);
  nor NOR2_23(g3927,g3382,g3383);
  nor NOR2_24(g3903,g3505,g471);
  nor NOR2_25(g1418,g486,g943);
  nor NOR2_26(g4578,g4234,g3928);
  nor NOR2_27(g4261,g3762,g3295);
  nor NOR4_6(g6358,I8126,I8127,I8128,I8129);
  nor NOR2_28(g4589,g4180,g4183);
  nor NOR2_29(g1474,g760,g754);
  nor NOR2_30(g3956,g3337,g3349);
  nor NOR2_31(g4774,g4442,g4445);
  nor NOR2_32(g5091,g4698,g4701);
  nor NOR2_33(g4950,g1472,g4680);
  nor NOR2_34(g5227,g5019,g3559);
  nor NOR2_35(g4585,g4171,g4177);
  nor NOR2_36(g6494,g952,g6348);
  nor NOR3_2(g5048,g4819,g3491,g3559);
  nor NOR3_3(g3664,g2804,g2791,g2780);
  nor NOR2_37(g4000,g1250,g3425);
  nor NOR2_38(g5418,g5162,g5169);
  nor NOR2_39(g5093,g4683,g4684);
  nor NOR2_40(g4779,g4461,g4464);
  nor NOR2_41(g6492,g6348,g1734);
  nor NOR3_4(g4240,g1589,g1879,g3793);
  nor NOR2_42(g4596,g4184,g4186);
  nor NOR2_43(g1603,g1039,g658);
  nor NOR3_5(g2908,g536,g2010,g541);
  nor NOR2_44(g4581,g4156,g4160);
  nor NOR2_45(g5423,g5170,g5175);
  nor NOR2_46(g4432,g923,g4253);
  nor NOR4_7(g6436,g6385,g3733,g4328,g4080);
  nor NOR2_47(g4568,g4233,g3924);
  nor NOR4_8(g6335,I8079,I8080,I8081,I8082);
  nor NOR2_48(g5753,g1477,g5688);
  nor NOR2_49(g6495,g6354,g1775);
  nor NOR4_9(g6442,g6376,g4323,g4074,g4302);
  nor NOR4_10(g6429,g6376,g4086,g4074,g4302);
  nor NOR4_11(g6281,I7987,I7988,I7989,I7990);
  nor NOR4_12(g6449,g6385,g4334,g4328,g4080);
  nor NOR2_50(g4590,g4169,g4172);
  nor NOR2_51(g4877,g952,g4680);
  nor NOR4_13(g6445,g6376,g4323,g4309,g4068);
  nor NOR4_14(g5561,g5391,g1589,g3793,g1880);
  nor NOR2_52(g3929,g3373,g3376);
  nor NOR3_6(g1473,g944,g941,g939);
  nor NOR2_53(g4967,g4674,g952);
  nor NOR4_15(g6430,g6385,g3733,g4092,g4080);
  nor NOR2_54(g4993,g4674,g1477);
  nor NOR4_16(g6448,g6376,g4323,g4309,g4302);
  nor NOR3_7(g3647,g2731,g2719,g2698);
  nor NOR2_55(g3925,g3303,g3315);
  nor NOR2_56(g5731,g952,g5688);
  nor NOR2_57(g3959,g3352,g3360);
  nor NOR2_58(g1481,g815,g809);
  nor NOR3_8(g3656,g2769,g2757,g2745);
  nor NOR2_59(g4245,g3759,g3288);
  nor NOR2_60(g3930,g3317,g3328);
  nor NOR2_61(g5249,g4868,g4870);
  nor NOR2_62(g3966,g3329,g3339);
  nor NOR4_17(g6400,I8208,I8209,I8210,I8211);
  nor NOR2_63(g4266,g3757,g3283);
  nor NOR4_18(g6451,g6385,g4334,g4328,g4314);
  nor NOR3_9(g5324,g5069,g4410,g766);
  nor NOR4_19(g6443,g6385,g4334,g4092,g4080);
  nor NOR2_64(g5088,g4691,g4697);
  nor NOR2_65(g3958,g3316,g3326);
  nor NOR2_66(g4241,g3774,g3341);
  nor NOR4_20(g6432,g6376,g4086,g4309,g4068);
  nor NOR4_21(g6357,I8117,I8118,I8119,I8120);
  nor NOR2_67(g3923,g3378,g3381);
  nor NOR2_68(g6075,g269,g5863);
  nor NOR2_69(g3934,g3377,g3379);
  nor NOR4_22(g6439,g6385,g3733,g4328,g4314);
  nor NOR2_70(g4272,g3767,g3319);
  nor NOR2_71(g1879,g1603,g1416);
  nor NOR3_10(g5325,g5077,g4416,g821);
  nor NOR4_23(g6435,g6376,g4086,g4309,g4302);
  nor NOR2_72(g4586,g4161,g4165);
  nor NOR2_73(g3939,g3340,g3351);
  nor NOR4_24(g6438,g6376,g4323,g4074,g4068);
  nor NOR2_74(g1518,g980,g965);
  nor NOR2_75(g4239,g3763,g3296);
  nor NOR2_76(g4591,g4178,g4181);

endmodule
